/*  Concrete parameterizations of argmin for testing.
 * 
 *  Copyright (c) 2016, Stephen Longfield, stephenlongfield.com
 * 
 *  This program is free software: you can redistribute it and/or modify
 *  it under the terms of the GNU General Public License as published by
 *  the Free Software Foundation, either version 3 of the License, or
 *  (at your option) any later version.
 *
 *  This program is distributed in the hope that it will be useful,
 *  but WITHOUT ANY WARRANTY; without even the implied warranty of
 *  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *  GNU General Public License for more details.
 *
 *  You should have received a copy of the GNU General Public License
 *  along with this program.  If not, see <http://www.gnu.org/licenses/>.
 *
 */

`include "argmin_10.v"

module argmin_test(
  input clk,
  input rst,
  input wire  [10*32-1:0] inp,
  output wire [31:0] outp,
  output wire [3:0] outp_addr
  );

  argmin_10#(.WIDTH(32)) am(clk, rst, inp, outp, outp_addr);

endmodule
