// Combinatorial MinDistance 
// 
// Generater written by: 
// Stephen Longfield, Dec 15, 2008 
// Generated fresh on 2009-01-23

module mindistance4(clk, reset, lham, rham, dout); 

  parameter HAMMING_TOTAL_SIZE =3599;
  parameter HAMMING_DEPTH = 11;
  parameter MAX_DISPARITY = 89;
  parameter DISPARITY_DEPTH = 6;
		
	
  input clk;
  input reset;
  input [HAMMING_TOTAL_SIZE:0] lham;
  input [HAMMING_TOTAL_SIZE:0] rham;
  output reg [DISPARITY_DEPTH:0] dout;

  reg [HAMMING_TOTAL_SIZE:0] rham_shift [MAX_DISPARITY:0];
  wire [HAMMING_DEPTH:0] distances [MAX_DISPARITY:0];


  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts0 (clk,reset,lham^rham_shift[0],distances[0]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts1 (clk,reset,lham^rham_shift[1],distances[1]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts2 (clk,reset,lham^rham_shift[2],distances[2]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts3 (clk,reset,lham^rham_shift[3],distances[3]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts4 (clk,reset,lham^rham_shift[4],distances[4]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts5 (clk,reset,lham^rham_shift[5],distances[5]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts6 (clk,reset,lham^rham_shift[6],distances[6]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts7 (clk,reset,lham^rham_shift[7],distances[7]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts8 (clk,reset,lham^rham_shift[8],distances[8]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts9 (clk,reset,lham^rham_shift[9],distances[9]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts10 (clk,reset,lham^rham_shift[10],distances[10]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts11 (clk,reset,lham^rham_shift[11],distances[11]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts12 (clk,reset,lham^rham_shift[12],distances[12]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts13 (clk,reset,lham^rham_shift[13],distances[13]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts14 (clk,reset,lham^rham_shift[14],distances[14]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts15 (clk,reset,lham^rham_shift[15],distances[15]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts16 (clk,reset,lham^rham_shift[16],distances[16]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts17 (clk,reset,lham^rham_shift[17],distances[17]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts18 (clk,reset,lham^rham_shift[18],distances[18]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts19 (clk,reset,lham^rham_shift[19],distances[19]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts20 (clk,reset,lham^rham_shift[20],distances[20]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts21 (clk,reset,lham^rham_shift[21],distances[21]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts22 (clk,reset,lham^rham_shift[22],distances[22]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts23 (clk,reset,lham^rham_shift[23],distances[23]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts24 (clk,reset,lham^rham_shift[24],distances[24]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts25 (clk,reset,lham^rham_shift[25],distances[25]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts26 (clk,reset,lham^rham_shift[26],distances[26]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts27 (clk,reset,lham^rham_shift[27],distances[27]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts28 (clk,reset,lham^rham_shift[28],distances[28]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts29 (clk,reset,lham^rham_shift[29],distances[29]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts30 (clk,reset,lham^rham_shift[30],distances[30]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts31 (clk,reset,lham^rham_shift[31],distances[31]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts32 (clk,reset,lham^rham_shift[32],distances[32]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts33 (clk,reset,lham^rham_shift[33],distances[33]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts34 (clk,reset,lham^rham_shift[34],distances[34]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts35 (clk,reset,lham^rham_shift[35],distances[35]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts36 (clk,reset,lham^rham_shift[36],distances[36]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts37 (clk,reset,lham^rham_shift[37],distances[37]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts38 (clk,reset,lham^rham_shift[38],distances[38]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts39 (clk,reset,lham^rham_shift[39],distances[39]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts40 (clk,reset,lham^rham_shift[40],distances[40]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts41 (clk,reset,lham^rham_shift[41],distances[41]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts42 (clk,reset,lham^rham_shift[42],distances[42]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts43 (clk,reset,lham^rham_shift[43],distances[43]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts44 (clk,reset,lham^rham_shift[44],distances[44]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts45 (clk,reset,lham^rham_shift[45],distances[45]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts46 (clk,reset,lham^rham_shift[46],distances[46]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts47 (clk,reset,lham^rham_shift[47],distances[47]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts48 (clk,reset,lham^rham_shift[48],distances[48]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts49 (clk,reset,lham^rham_shift[49],distances[49]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts50 (clk,reset,lham^rham_shift[50],distances[50]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts51 (clk,reset,lham^rham_shift[51],distances[51]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts52 (clk,reset,lham^rham_shift[52],distances[52]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts53 (clk,reset,lham^rham_shift[53],distances[53]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts54 (clk,reset,lham^rham_shift[54],distances[54]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts55 (clk,reset,lham^rham_shift[55],distances[55]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts56 (clk,reset,lham^rham_shift[56],distances[56]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts57 (clk,reset,lham^rham_shift[57],distances[57]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts58 (clk,reset,lham^rham_shift[58],distances[58]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts59 (clk,reset,lham^rham_shift[59],distances[59]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts60 (clk,reset,lham^rham_shift[60],distances[60]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts61 (clk,reset,lham^rham_shift[61],distances[61]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts62 (clk,reset,lham^rham_shift[62],distances[62]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts63 (clk,reset,lham^rham_shift[63],distances[63]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts64 (clk,reset,lham^rham_shift[64],distances[64]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts65 (clk,reset,lham^rham_shift[65],distances[65]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts66 (clk,reset,lham^rham_shift[66],distances[66]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts67 (clk,reset,lham^rham_shift[67],distances[67]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts68 (clk,reset,lham^rham_shift[68],distances[68]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts69 (clk,reset,lham^rham_shift[69],distances[69]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts70 (clk,reset,lham^rham_shift[70],distances[70]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts71 (clk,reset,lham^rham_shift[71],distances[71]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts72 (clk,reset,lham^rham_shift[72],distances[72]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts73 (clk,reset,lham^rham_shift[73],distances[73]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts74 (clk,reset,lham^rham_shift[74],distances[74]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts75 (clk,reset,lham^rham_shift[75],distances[75]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts76 (clk,reset,lham^rham_shift[76],distances[76]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts77 (clk,reset,lham^rham_shift[77],distances[77]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts78 (clk,reset,lham^rham_shift[78],distances[78]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts79 (clk,reset,lham^rham_shift[79],distances[79]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts80 (clk,reset,lham^rham_shift[80],distances[80]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts81 (clk,reset,lham^rham_shift[81],distances[81]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts82 (clk,reset,lham^rham_shift[82],distances[82]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts83 (clk,reset,lham^rham_shift[83],distances[83]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts84 (clk,reset,lham^rham_shift[84],distances[84]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts85 (clk,reset,lham^rham_shift[85],distances[85]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts86 (clk,reset,lham^rham_shift[86],distances[86]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts87 (clk,reset,lham^rham_shift[87],distances[87]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts88 (clk,reset,lham^rham_shift[88],distances[88]);

  treesum #(.HAMMING_TOTAL_SIZE(HAMMING_TOTAL_SIZE), .HAMMING_DEPTH(HAMMING_DEPTH))
                    ts89 (clk,reset,lham^rham_shift[89],distances[89]);

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      dout <= 0;

      rham_shift[0] <= 0;
      rham_shift[1] <= 0;
      rham_shift[2] <= 0;
      rham_shift[3] <= 0;
      rham_shift[4] <= 0;
      rham_shift[5] <= 0;
      rham_shift[6] <= 0;
      rham_shift[7] <= 0;
      rham_shift[8] <= 0;
      rham_shift[9] <= 0;
      rham_shift[10] <= 0;
      rham_shift[11] <= 0;
      rham_shift[12] <= 0;
      rham_shift[13] <= 0;
      rham_shift[14] <= 0;
      rham_shift[15] <= 0;
      rham_shift[16] <= 0;
      rham_shift[17] <= 0;
      rham_shift[18] <= 0;
      rham_shift[19] <= 0;
      rham_shift[20] <= 0;
      rham_shift[21] <= 0;
      rham_shift[22] <= 0;
      rham_shift[23] <= 0;
      rham_shift[24] <= 0;
      rham_shift[25] <= 0;
      rham_shift[26] <= 0;
      rham_shift[27] <= 0;
      rham_shift[28] <= 0;
      rham_shift[29] <= 0;
      rham_shift[30] <= 0;
      rham_shift[31] <= 0;
      rham_shift[32] <= 0;
      rham_shift[33] <= 0;
      rham_shift[34] <= 0;
      rham_shift[35] <= 0;
      rham_shift[36] <= 0;
      rham_shift[37] <= 0;
      rham_shift[38] <= 0;
      rham_shift[39] <= 0;
      rham_shift[40] <= 0;
      rham_shift[41] <= 0;
      rham_shift[42] <= 0;
      rham_shift[43] <= 0;
      rham_shift[44] <= 0;
      rham_shift[45] <= 0;
      rham_shift[46] <= 0;
      rham_shift[47] <= 0;
      rham_shift[48] <= 0;
      rham_shift[49] <= 0;
      rham_shift[50] <= 0;
      rham_shift[51] <= 0;
      rham_shift[52] <= 0;
      rham_shift[53] <= 0;
      rham_shift[54] <= 0;
      rham_shift[55] <= 0;
      rham_shift[56] <= 0;
      rham_shift[57] <= 0;
      rham_shift[58] <= 0;
      rham_shift[59] <= 0;
      rham_shift[60] <= 0;
      rham_shift[61] <= 0;
      rham_shift[62] <= 0;
      rham_shift[63] <= 0;
      rham_shift[64] <= 0;
      rham_shift[65] <= 0;
      rham_shift[66] <= 0;
      rham_shift[67] <= 0;
      rham_shift[68] <= 0;
      rham_shift[69] <= 0;
      rham_shift[70] <= 0;
      rham_shift[71] <= 0;
      rham_shift[72] <= 0;
      rham_shift[73] <= 0;
      rham_shift[74] <= 0;
      rham_shift[75] <= 0;
      rham_shift[76] <= 0;
      rham_shift[77] <= 0;
      rham_shift[78] <= 0;
      rham_shift[79] <= 0;
      rham_shift[80] <= 0;
      rham_shift[81] <= 0;
      rham_shift[82] <= 0;
      rham_shift[83] <= 0;
      rham_shift[84] <= 0;
      rham_shift[85] <= 0;
      rham_shift[86] <= 0;
      rham_shift[87] <= 0;
      rham_shift[88] <= 0;
      rham_shift[89] <= 0;
    end else begin
      rham_shift[0] <= rham;
      rham_shift[1] <= rham_shift[0];
      rham_shift[2] <= rham_shift[1];
      rham_shift[3] <= rham_shift[2];
      rham_shift[4] <= rham_shift[3];
      rham_shift[5] <= rham_shift[4];
      rham_shift[6] <= rham_shift[5];
      rham_shift[7] <= rham_shift[6];
      rham_shift[8] <= rham_shift[7];
      rham_shift[9] <= rham_shift[8];
      rham_shift[10] <= rham_shift[9];
      rham_shift[11] <= rham_shift[10];
      rham_shift[12] <= rham_shift[11];
      rham_shift[13] <= rham_shift[12];
      rham_shift[14] <= rham_shift[13];
      rham_shift[15] <= rham_shift[14];
      rham_shift[16] <= rham_shift[15];
      rham_shift[17] <= rham_shift[16];
      rham_shift[18] <= rham_shift[17];
      rham_shift[19] <= rham_shift[18];
      rham_shift[20] <= rham_shift[19];
      rham_shift[21] <= rham_shift[20];
      rham_shift[22] <= rham_shift[21];
      rham_shift[23] <= rham_shift[22];
      rham_shift[24] <= rham_shift[23];
      rham_shift[25] <= rham_shift[24];
      rham_shift[26] <= rham_shift[25];
      rham_shift[27] <= rham_shift[26];
      rham_shift[28] <= rham_shift[27];
      rham_shift[29] <= rham_shift[28];
      rham_shift[30] <= rham_shift[29];
      rham_shift[31] <= rham_shift[30];
      rham_shift[32] <= rham_shift[31];
      rham_shift[33] <= rham_shift[32];
      rham_shift[34] <= rham_shift[33];
      rham_shift[35] <= rham_shift[34];
      rham_shift[36] <= rham_shift[35];
      rham_shift[37] <= rham_shift[36];
      rham_shift[38] <= rham_shift[37];
      rham_shift[39] <= rham_shift[38];
      rham_shift[40] <= rham_shift[39];
      rham_shift[41] <= rham_shift[40];
      rham_shift[42] <= rham_shift[41];
      rham_shift[43] <= rham_shift[42];
      rham_shift[44] <= rham_shift[43];
      rham_shift[45] <= rham_shift[44];
      rham_shift[46] <= rham_shift[45];
      rham_shift[47] <= rham_shift[46];
      rham_shift[48] <= rham_shift[47];
      rham_shift[49] <= rham_shift[48];
      rham_shift[50] <= rham_shift[49];
      rham_shift[51] <= rham_shift[50];
      rham_shift[52] <= rham_shift[51];
      rham_shift[53] <= rham_shift[52];
      rham_shift[54] <= rham_shift[53];
      rham_shift[55] <= rham_shift[54];
      rham_shift[56] <= rham_shift[55];
      rham_shift[57] <= rham_shift[56];
      rham_shift[58] <= rham_shift[57];
      rham_shift[59] <= rham_shift[58];
      rham_shift[60] <= rham_shift[59];
      rham_shift[61] <= rham_shift[60];
      rham_shift[62] <= rham_shift[61];
      rham_shift[63] <= rham_shift[62];
      rham_shift[64] <= rham_shift[63];
      rham_shift[65] <= rham_shift[64];
      rham_shift[66] <= rham_shift[65];
      rham_shift[67] <= rham_shift[66];
      rham_shift[68] <= rham_shift[67];
      rham_shift[69] <= rham_shift[68];
      rham_shift[70] <= rham_shift[69];
      rham_shift[71] <= rham_shift[70];
      rham_shift[72] <= rham_shift[71];
      rham_shift[73] <= rham_shift[72];
      rham_shift[74] <= rham_shift[73];
      rham_shift[75] <= rham_shift[74];
      rham_shift[76] <= rham_shift[75];
      rham_shift[77] <= rham_shift[76];
      rham_shift[78] <= rham_shift[77];
      rham_shift[79] <= rham_shift[78];
      rham_shift[80] <= rham_shift[79];
      rham_shift[81] <= rham_shift[80];
      rham_shift[82] <= rham_shift[81];
      rham_shift[83] <= rham_shift[82];
      rham_shift[84] <= rham_shift[83];
      rham_shift[85] <= rham_shift[84];
      rham_shift[86] <= rham_shift[85];
      rham_shift[87] <= rham_shift[86];
      rham_shift[88] <= rham_shift[87];
      rham_shift[89] <= rham_shift[88];

      if ((distances[0] < distances[1]) && (distances[0] < distances[2]) && (distances[0] < distances[3]) && (distances[0] < distances[4]) && (distances[0] < distances[5]) && (distances[0] < distances[6]) && (distances[0] < distances[7]) && (distances[0] < distances[8]) && (distances[0] < distances[9]) && (distances[0] < distances[10]) && (distances[0] < distances[11]) && (distances[0] < distances[12]) && (distances[0] < distances[13]) && (distances[0] < distances[14]) && (distances[0] < distances[15]) && (distances[0] < distances[16]) && (distances[0] < distances[17]) && (distances[0] < distances[18]) && (distances[0] < distances[19]) && (distances[0] < distances[20]) && (distances[0] < distances[21]) && (distances[0] < distances[22]) && (distances[0] < distances[23]) && (distances[0] < distances[24]) && (distances[0] < distances[25]) && (distances[0] < distances[26]) && (distances[0] < distances[27]) && (distances[0] < distances[28]) && (distances[0] < distances[29]) && (distances[0] < distances[30]) && (distances[0] < distances[31]) && (distances[0] < distances[32]) && (distances[0] < distances[33]) && (distances[0] < distances[34]) && (distances[0] < distances[35]) && (distances[0] < distances[36]) && (distances[0] < distances[37]) && (distances[0] < distances[38]) && (distances[0] < distances[39]) && (distances[0] < distances[40]) && (distances[0] < distances[41]) && (distances[0] < distances[42]) && (distances[0] < distances[43]) && (distances[0] < distances[44]) && (distances[0] < distances[45]) && (distances[0] < distances[46]) && (distances[0] < distances[47]) && (distances[0] < distances[48]) && (distances[0] < distances[49]) && (distances[0] < distances[50]) && (distances[0] < distances[51]) && (distances[0] < distances[52]) && (distances[0] < distances[53]) && (distances[0] < distances[54]) && (distances[0] < distances[55]) && (distances[0] < distances[56]) && (distances[0] < distances[57]) && (distances[0] < distances[58]) && (distances[0] < distances[59]) && (distances[0] < distances[60]) && (distances[0] < distances[61]) && (distances[0] < distances[62]) && (distances[0] < distances[63]) && (distances[0] < distances[64]) && (distances[0] < distances[65]) && (distances[0] < distances[66]) && (distances[0] < distances[67]) && (distances[0] < distances[68]) && (distances[0] < distances[69]) && (distances[0] < distances[70]) && (distances[0] < distances[71]) && (distances[0] < distances[72]) && (distances[0] < distances[73]) && (distances[0] < distances[74]) && (distances[0] < distances[75]) && (distances[0] < distances[76]) && (distances[0] < distances[77]) && (distances[0] < distances[78]) && (distances[0] < distances[79]) && (distances[0] < distances[80]) && (distances[0] < distances[81]) && (distances[0] < distances[82]) && (distances[0] < distances[83]) && (distances[0] < distances[84]) && (distances[0] < distances[85]) && (distances[0] < distances[86]) && (distances[0] < distances[87]) && (distances[0] < distances[88]) && (distances[0] < distances[89])) begin
        dout <= 0;
      end else if((distances[1] < distances[2]) && (distances[1] < distances[3]) && (distances[1] < distances[4]) && (distances[1] < distances[5]) && (distances[1] < distances[6]) && (distances[1] < distances[7]) && (distances[1] < distances[8]) && (distances[1] < distances[9]) && (distances[1] < distances[10]) && (distances[1] < distances[11]) && (distances[1] < distances[12]) && (distances[1] < distances[13]) && (distances[1] < distances[14]) && (distances[1] < distances[15]) && (distances[1] < distances[16]) && (distances[1] < distances[17]) && (distances[1] < distances[18]) && (distances[1] < distances[19]) && (distances[1] < distances[20]) && (distances[1] < distances[21]) && (distances[1] < distances[22]) && (distances[1] < distances[23]) && (distances[1] < distances[24]) && (distances[1] < distances[25]) && (distances[1] < distances[26]) && (distances[1] < distances[27]) && (distances[1] < distances[28]) && (distances[1] < distances[29]) && (distances[1] < distances[30]) && (distances[1] < distances[31]) && (distances[1] < distances[32]) && (distances[1] < distances[33]) && (distances[1] < distances[34]) && (distances[1] < distances[35]) && (distances[1] < distances[36]) && (distances[1] < distances[37]) && (distances[1] < distances[38]) && (distances[1] < distances[39]) && (distances[1] < distances[40]) && (distances[1] < distances[41]) && (distances[1] < distances[42]) && (distances[1] < distances[43]) && (distances[1] < distances[44]) && (distances[1] < distances[45]) && (distances[1] < distances[46]) && (distances[1] < distances[47]) && (distances[1] < distances[48]) && (distances[1] < distances[49]) && (distances[1] < distances[50]) && (distances[1] < distances[51]) && (distances[1] < distances[52]) && (distances[1] < distances[53]) && (distances[1] < distances[54]) && (distances[1] < distances[55]) && (distances[1] < distances[56]) && (distances[1] < distances[57]) && (distances[1] < distances[58]) && (distances[1] < distances[59]) && (distances[1] < distances[60]) && (distances[1] < distances[61]) && (distances[1] < distances[62]) && (distances[1] < distances[63]) && (distances[1] < distances[64]) && (distances[1] < distances[65]) && (distances[1] < distances[66]) && (distances[1] < distances[67]) && (distances[1] < distances[68]) && (distances[1] < distances[69]) && (distances[1] < distances[70]) && (distances[1] < distances[71]) && (distances[1] < distances[72]) && (distances[1] < distances[73]) && (distances[1] < distances[74]) && (distances[1] < distances[75]) && (distances[1] < distances[76]) && (distances[1] < distances[77]) && (distances[1] < distances[78]) && (distances[1] < distances[79]) && (distances[1] < distances[80]) && (distances[1] < distances[81]) && (distances[1] < distances[82]) && (distances[1] < distances[83]) && (distances[1] < distances[84]) && (distances[1] < distances[85]) && (distances[1] < distances[86]) && (distances[1] < distances[87]) && (distances[1] < distances[88]) && (distances[1] < distances[89])) begin
        dout <= 1;
      end else if((distances[2] < distances[3]) && (distances[2] < distances[4]) && (distances[2] < distances[5]) && (distances[2] < distances[6]) && (distances[2] < distances[7]) && (distances[2] < distances[8]) && (distances[2] < distances[9]) && (distances[2] < distances[10]) && (distances[2] < distances[11]) && (distances[2] < distances[12]) && (distances[2] < distances[13]) && (distances[2] < distances[14]) && (distances[2] < distances[15]) && (distances[2] < distances[16]) && (distances[2] < distances[17]) && (distances[2] < distances[18]) && (distances[2] < distances[19]) && (distances[2] < distances[20]) && (distances[2] < distances[21]) && (distances[2] < distances[22]) && (distances[2] < distances[23]) && (distances[2] < distances[24]) && (distances[2] < distances[25]) && (distances[2] < distances[26]) && (distances[2] < distances[27]) && (distances[2] < distances[28]) && (distances[2] < distances[29]) && (distances[2] < distances[30]) && (distances[2] < distances[31]) && (distances[2] < distances[32]) && (distances[2] < distances[33]) && (distances[2] < distances[34]) && (distances[2] < distances[35]) && (distances[2] < distances[36]) && (distances[2] < distances[37]) && (distances[2] < distances[38]) && (distances[2] < distances[39]) && (distances[2] < distances[40]) && (distances[2] < distances[41]) && (distances[2] < distances[42]) && (distances[2] < distances[43]) && (distances[2] < distances[44]) && (distances[2] < distances[45]) && (distances[2] < distances[46]) && (distances[2] < distances[47]) && (distances[2] < distances[48]) && (distances[2] < distances[49]) && (distances[2] < distances[50]) && (distances[2] < distances[51]) && (distances[2] < distances[52]) && (distances[2] < distances[53]) && (distances[2] < distances[54]) && (distances[2] < distances[55]) && (distances[2] < distances[56]) && (distances[2] < distances[57]) && (distances[2] < distances[58]) && (distances[2] < distances[59]) && (distances[2] < distances[60]) && (distances[2] < distances[61]) && (distances[2] < distances[62]) && (distances[2] < distances[63]) && (distances[2] < distances[64]) && (distances[2] < distances[65]) && (distances[2] < distances[66]) && (distances[2] < distances[67]) && (distances[2] < distances[68]) && (distances[2] < distances[69]) && (distances[2] < distances[70]) && (distances[2] < distances[71]) && (distances[2] < distances[72]) && (distances[2] < distances[73]) && (distances[2] < distances[74]) && (distances[2] < distances[75]) && (distances[2] < distances[76]) && (distances[2] < distances[77]) && (distances[2] < distances[78]) && (distances[2] < distances[79]) && (distances[2] < distances[80]) && (distances[2] < distances[81]) && (distances[2] < distances[82]) && (distances[2] < distances[83]) && (distances[2] < distances[84]) && (distances[2] < distances[85]) && (distances[2] < distances[86]) && (distances[2] < distances[87]) && (distances[2] < distances[88]) && (distances[2] < distances[89])) begin
        dout <= 2;
      end else if((distances[3] < distances[4]) && (distances[3] < distances[5]) && (distances[3] < distances[6]) && (distances[3] < distances[7]) && (distances[3] < distances[8]) && (distances[3] < distances[9]) && (distances[3] < distances[10]) && (distances[3] < distances[11]) && (distances[3] < distances[12]) && (distances[3] < distances[13]) && (distances[3] < distances[14]) && (distances[3] < distances[15]) && (distances[3] < distances[16]) && (distances[3] < distances[17]) && (distances[3] < distances[18]) && (distances[3] < distances[19]) && (distances[3] < distances[20]) && (distances[3] < distances[21]) && (distances[3] < distances[22]) && (distances[3] < distances[23]) && (distances[3] < distances[24]) && (distances[3] < distances[25]) && (distances[3] < distances[26]) && (distances[3] < distances[27]) && (distances[3] < distances[28]) && (distances[3] < distances[29]) && (distances[3] < distances[30]) && (distances[3] < distances[31]) && (distances[3] < distances[32]) && (distances[3] < distances[33]) && (distances[3] < distances[34]) && (distances[3] < distances[35]) && (distances[3] < distances[36]) && (distances[3] < distances[37]) && (distances[3] < distances[38]) && (distances[3] < distances[39]) && (distances[3] < distances[40]) && (distances[3] < distances[41]) && (distances[3] < distances[42]) && (distances[3] < distances[43]) && (distances[3] < distances[44]) && (distances[3] < distances[45]) && (distances[3] < distances[46]) && (distances[3] < distances[47]) && (distances[3] < distances[48]) && (distances[3] < distances[49]) && (distances[3] < distances[50]) && (distances[3] < distances[51]) && (distances[3] < distances[52]) && (distances[3] < distances[53]) && (distances[3] < distances[54]) && (distances[3] < distances[55]) && (distances[3] < distances[56]) && (distances[3] < distances[57]) && (distances[3] < distances[58]) && (distances[3] < distances[59]) && (distances[3] < distances[60]) && (distances[3] < distances[61]) && (distances[3] < distances[62]) && (distances[3] < distances[63]) && (distances[3] < distances[64]) && (distances[3] < distances[65]) && (distances[3] < distances[66]) && (distances[3] < distances[67]) && (distances[3] < distances[68]) && (distances[3] < distances[69]) && (distances[3] < distances[70]) && (distances[3] < distances[71]) && (distances[3] < distances[72]) && (distances[3] < distances[73]) && (distances[3] < distances[74]) && (distances[3] < distances[75]) && (distances[3] < distances[76]) && (distances[3] < distances[77]) && (distances[3] < distances[78]) && (distances[3] < distances[79]) && (distances[3] < distances[80]) && (distances[3] < distances[81]) && (distances[3] < distances[82]) && (distances[3] < distances[83]) && (distances[3] < distances[84]) && (distances[3] < distances[85]) && (distances[3] < distances[86]) && (distances[3] < distances[87]) && (distances[3] < distances[88]) && (distances[3] < distances[89])) begin
        dout <= 3;
      end else if((distances[4] < distances[5]) && (distances[4] < distances[6]) && (distances[4] < distances[7]) && (distances[4] < distances[8]) && (distances[4] < distances[9]) && (distances[4] < distances[10]) && (distances[4] < distances[11]) && (distances[4] < distances[12]) && (distances[4] < distances[13]) && (distances[4] < distances[14]) && (distances[4] < distances[15]) && (distances[4] < distances[16]) && (distances[4] < distances[17]) && (distances[4] < distances[18]) && (distances[4] < distances[19]) && (distances[4] < distances[20]) && (distances[4] < distances[21]) && (distances[4] < distances[22]) && (distances[4] < distances[23]) && (distances[4] < distances[24]) && (distances[4] < distances[25]) && (distances[4] < distances[26]) && (distances[4] < distances[27]) && (distances[4] < distances[28]) && (distances[4] < distances[29]) && (distances[4] < distances[30]) && (distances[4] < distances[31]) && (distances[4] < distances[32]) && (distances[4] < distances[33]) && (distances[4] < distances[34]) && (distances[4] < distances[35]) && (distances[4] < distances[36]) && (distances[4] < distances[37]) && (distances[4] < distances[38]) && (distances[4] < distances[39]) && (distances[4] < distances[40]) && (distances[4] < distances[41]) && (distances[4] < distances[42]) && (distances[4] < distances[43]) && (distances[4] < distances[44]) && (distances[4] < distances[45]) && (distances[4] < distances[46]) && (distances[4] < distances[47]) && (distances[4] < distances[48]) && (distances[4] < distances[49]) && (distances[4] < distances[50]) && (distances[4] < distances[51]) && (distances[4] < distances[52]) && (distances[4] < distances[53]) && (distances[4] < distances[54]) && (distances[4] < distances[55]) && (distances[4] < distances[56]) && (distances[4] < distances[57]) && (distances[4] < distances[58]) && (distances[4] < distances[59]) && (distances[4] < distances[60]) && (distances[4] < distances[61]) && (distances[4] < distances[62]) && (distances[4] < distances[63]) && (distances[4] < distances[64]) && (distances[4] < distances[65]) && (distances[4] < distances[66]) && (distances[4] < distances[67]) && (distances[4] < distances[68]) && (distances[4] < distances[69]) && (distances[4] < distances[70]) && (distances[4] < distances[71]) && (distances[4] < distances[72]) && (distances[4] < distances[73]) && (distances[4] < distances[74]) && (distances[4] < distances[75]) && (distances[4] < distances[76]) && (distances[4] < distances[77]) && (distances[4] < distances[78]) && (distances[4] < distances[79]) && (distances[4] < distances[80]) && (distances[4] < distances[81]) && (distances[4] < distances[82]) && (distances[4] < distances[83]) && (distances[4] < distances[84]) && (distances[4] < distances[85]) && (distances[4] < distances[86]) && (distances[4] < distances[87]) && (distances[4] < distances[88]) && (distances[4] < distances[89])) begin
        dout <= 4;
      end else if((distances[5] < distances[6]) && (distances[5] < distances[7]) && (distances[5] < distances[8]) && (distances[5] < distances[9]) && (distances[5] < distances[10]) && (distances[5] < distances[11]) && (distances[5] < distances[12]) && (distances[5] < distances[13]) && (distances[5] < distances[14]) && (distances[5] < distances[15]) && (distances[5] < distances[16]) && (distances[5] < distances[17]) && (distances[5] < distances[18]) && (distances[5] < distances[19]) && (distances[5] < distances[20]) && (distances[5] < distances[21]) && (distances[5] < distances[22]) && (distances[5] < distances[23]) && (distances[5] < distances[24]) && (distances[5] < distances[25]) && (distances[5] < distances[26]) && (distances[5] < distances[27]) && (distances[5] < distances[28]) && (distances[5] < distances[29]) && (distances[5] < distances[30]) && (distances[5] < distances[31]) && (distances[5] < distances[32]) && (distances[5] < distances[33]) && (distances[5] < distances[34]) && (distances[5] < distances[35]) && (distances[5] < distances[36]) && (distances[5] < distances[37]) && (distances[5] < distances[38]) && (distances[5] < distances[39]) && (distances[5] < distances[40]) && (distances[5] < distances[41]) && (distances[5] < distances[42]) && (distances[5] < distances[43]) && (distances[5] < distances[44]) && (distances[5] < distances[45]) && (distances[5] < distances[46]) && (distances[5] < distances[47]) && (distances[5] < distances[48]) && (distances[5] < distances[49]) && (distances[5] < distances[50]) && (distances[5] < distances[51]) && (distances[5] < distances[52]) && (distances[5] < distances[53]) && (distances[5] < distances[54]) && (distances[5] < distances[55]) && (distances[5] < distances[56]) && (distances[5] < distances[57]) && (distances[5] < distances[58]) && (distances[5] < distances[59]) && (distances[5] < distances[60]) && (distances[5] < distances[61]) && (distances[5] < distances[62]) && (distances[5] < distances[63]) && (distances[5] < distances[64]) && (distances[5] < distances[65]) && (distances[5] < distances[66]) && (distances[5] < distances[67]) && (distances[5] < distances[68]) && (distances[5] < distances[69]) && (distances[5] < distances[70]) && (distances[5] < distances[71]) && (distances[5] < distances[72]) && (distances[5] < distances[73]) && (distances[5] < distances[74]) && (distances[5] < distances[75]) && (distances[5] < distances[76]) && (distances[5] < distances[77]) && (distances[5] < distances[78]) && (distances[5] < distances[79]) && (distances[5] < distances[80]) && (distances[5] < distances[81]) && (distances[5] < distances[82]) && (distances[5] < distances[83]) && (distances[5] < distances[84]) && (distances[5] < distances[85]) && (distances[5] < distances[86]) && (distances[5] < distances[87]) && (distances[5] < distances[88]) && (distances[5] < distances[89])) begin
        dout <= 5;
      end else if((distances[6] < distances[7]) && (distances[6] < distances[8]) && (distances[6] < distances[9]) && (distances[6] < distances[10]) && (distances[6] < distances[11]) && (distances[6] < distances[12]) && (distances[6] < distances[13]) && (distances[6] < distances[14]) && (distances[6] < distances[15]) && (distances[6] < distances[16]) && (distances[6] < distances[17]) && (distances[6] < distances[18]) && (distances[6] < distances[19]) && (distances[6] < distances[20]) && (distances[6] < distances[21]) && (distances[6] < distances[22]) && (distances[6] < distances[23]) && (distances[6] < distances[24]) && (distances[6] < distances[25]) && (distances[6] < distances[26]) && (distances[6] < distances[27]) && (distances[6] < distances[28]) && (distances[6] < distances[29]) && (distances[6] < distances[30]) && (distances[6] < distances[31]) && (distances[6] < distances[32]) && (distances[6] < distances[33]) && (distances[6] < distances[34]) && (distances[6] < distances[35]) && (distances[6] < distances[36]) && (distances[6] < distances[37]) && (distances[6] < distances[38]) && (distances[6] < distances[39]) && (distances[6] < distances[40]) && (distances[6] < distances[41]) && (distances[6] < distances[42]) && (distances[6] < distances[43]) && (distances[6] < distances[44]) && (distances[6] < distances[45]) && (distances[6] < distances[46]) && (distances[6] < distances[47]) && (distances[6] < distances[48]) && (distances[6] < distances[49]) && (distances[6] < distances[50]) && (distances[6] < distances[51]) && (distances[6] < distances[52]) && (distances[6] < distances[53]) && (distances[6] < distances[54]) && (distances[6] < distances[55]) && (distances[6] < distances[56]) && (distances[6] < distances[57]) && (distances[6] < distances[58]) && (distances[6] < distances[59]) && (distances[6] < distances[60]) && (distances[6] < distances[61]) && (distances[6] < distances[62]) && (distances[6] < distances[63]) && (distances[6] < distances[64]) && (distances[6] < distances[65]) && (distances[6] < distances[66]) && (distances[6] < distances[67]) && (distances[6] < distances[68]) && (distances[6] < distances[69]) && (distances[6] < distances[70]) && (distances[6] < distances[71]) && (distances[6] < distances[72]) && (distances[6] < distances[73]) && (distances[6] < distances[74]) && (distances[6] < distances[75]) && (distances[6] < distances[76]) && (distances[6] < distances[77]) && (distances[6] < distances[78]) && (distances[6] < distances[79]) && (distances[6] < distances[80]) && (distances[6] < distances[81]) && (distances[6] < distances[82]) && (distances[6] < distances[83]) && (distances[6] < distances[84]) && (distances[6] < distances[85]) && (distances[6] < distances[86]) && (distances[6] < distances[87]) && (distances[6] < distances[88]) && (distances[6] < distances[89])) begin
        dout <= 6;
      end else if((distances[7] < distances[8]) && (distances[7] < distances[9]) && (distances[7] < distances[10]) && (distances[7] < distances[11]) && (distances[7] < distances[12]) && (distances[7] < distances[13]) && (distances[7] < distances[14]) && (distances[7] < distances[15]) && (distances[7] < distances[16]) && (distances[7] < distances[17]) && (distances[7] < distances[18]) && (distances[7] < distances[19]) && (distances[7] < distances[20]) && (distances[7] < distances[21]) && (distances[7] < distances[22]) && (distances[7] < distances[23]) && (distances[7] < distances[24]) && (distances[7] < distances[25]) && (distances[7] < distances[26]) && (distances[7] < distances[27]) && (distances[7] < distances[28]) && (distances[7] < distances[29]) && (distances[7] < distances[30]) && (distances[7] < distances[31]) && (distances[7] < distances[32]) && (distances[7] < distances[33]) && (distances[7] < distances[34]) && (distances[7] < distances[35]) && (distances[7] < distances[36]) && (distances[7] < distances[37]) && (distances[7] < distances[38]) && (distances[7] < distances[39]) && (distances[7] < distances[40]) && (distances[7] < distances[41]) && (distances[7] < distances[42]) && (distances[7] < distances[43]) && (distances[7] < distances[44]) && (distances[7] < distances[45]) && (distances[7] < distances[46]) && (distances[7] < distances[47]) && (distances[7] < distances[48]) && (distances[7] < distances[49]) && (distances[7] < distances[50]) && (distances[7] < distances[51]) && (distances[7] < distances[52]) && (distances[7] < distances[53]) && (distances[7] < distances[54]) && (distances[7] < distances[55]) && (distances[7] < distances[56]) && (distances[7] < distances[57]) && (distances[7] < distances[58]) && (distances[7] < distances[59]) && (distances[7] < distances[60]) && (distances[7] < distances[61]) && (distances[7] < distances[62]) && (distances[7] < distances[63]) && (distances[7] < distances[64]) && (distances[7] < distances[65]) && (distances[7] < distances[66]) && (distances[7] < distances[67]) && (distances[7] < distances[68]) && (distances[7] < distances[69]) && (distances[7] < distances[70]) && (distances[7] < distances[71]) && (distances[7] < distances[72]) && (distances[7] < distances[73]) && (distances[7] < distances[74]) && (distances[7] < distances[75]) && (distances[7] < distances[76]) && (distances[7] < distances[77]) && (distances[7] < distances[78]) && (distances[7] < distances[79]) && (distances[7] < distances[80]) && (distances[7] < distances[81]) && (distances[7] < distances[82]) && (distances[7] < distances[83]) && (distances[7] < distances[84]) && (distances[7] < distances[85]) && (distances[7] < distances[86]) && (distances[7] < distances[87]) && (distances[7] < distances[88]) && (distances[7] < distances[89])) begin
        dout <= 7;
      end else if((distances[8] < distances[9]) && (distances[8] < distances[10]) && (distances[8] < distances[11]) && (distances[8] < distances[12]) && (distances[8] < distances[13]) && (distances[8] < distances[14]) && (distances[8] < distances[15]) && (distances[8] < distances[16]) && (distances[8] < distances[17]) && (distances[8] < distances[18]) && (distances[8] < distances[19]) && (distances[8] < distances[20]) && (distances[8] < distances[21]) && (distances[8] < distances[22]) && (distances[8] < distances[23]) && (distances[8] < distances[24]) && (distances[8] < distances[25]) && (distances[8] < distances[26]) && (distances[8] < distances[27]) && (distances[8] < distances[28]) && (distances[8] < distances[29]) && (distances[8] < distances[30]) && (distances[8] < distances[31]) && (distances[8] < distances[32]) && (distances[8] < distances[33]) && (distances[8] < distances[34]) && (distances[8] < distances[35]) && (distances[8] < distances[36]) && (distances[8] < distances[37]) && (distances[8] < distances[38]) && (distances[8] < distances[39]) && (distances[8] < distances[40]) && (distances[8] < distances[41]) && (distances[8] < distances[42]) && (distances[8] < distances[43]) && (distances[8] < distances[44]) && (distances[8] < distances[45]) && (distances[8] < distances[46]) && (distances[8] < distances[47]) && (distances[8] < distances[48]) && (distances[8] < distances[49]) && (distances[8] < distances[50]) && (distances[8] < distances[51]) && (distances[8] < distances[52]) && (distances[8] < distances[53]) && (distances[8] < distances[54]) && (distances[8] < distances[55]) && (distances[8] < distances[56]) && (distances[8] < distances[57]) && (distances[8] < distances[58]) && (distances[8] < distances[59]) && (distances[8] < distances[60]) && (distances[8] < distances[61]) && (distances[8] < distances[62]) && (distances[8] < distances[63]) && (distances[8] < distances[64]) && (distances[8] < distances[65]) && (distances[8] < distances[66]) && (distances[8] < distances[67]) && (distances[8] < distances[68]) && (distances[8] < distances[69]) && (distances[8] < distances[70]) && (distances[8] < distances[71]) && (distances[8] < distances[72]) && (distances[8] < distances[73]) && (distances[8] < distances[74]) && (distances[8] < distances[75]) && (distances[8] < distances[76]) && (distances[8] < distances[77]) && (distances[8] < distances[78]) && (distances[8] < distances[79]) && (distances[8] < distances[80]) && (distances[8] < distances[81]) && (distances[8] < distances[82]) && (distances[8] < distances[83]) && (distances[8] < distances[84]) && (distances[8] < distances[85]) && (distances[8] < distances[86]) && (distances[8] < distances[87]) && (distances[8] < distances[88]) && (distances[8] < distances[89])) begin
        dout <= 8;
      end else if((distances[9] < distances[10]) && (distances[9] < distances[11]) && (distances[9] < distances[12]) && (distances[9] < distances[13]) && (distances[9] < distances[14]) && (distances[9] < distances[15]) && (distances[9] < distances[16]) && (distances[9] < distances[17]) && (distances[9] < distances[18]) && (distances[9] < distances[19]) && (distances[9] < distances[20]) && (distances[9] < distances[21]) && (distances[9] < distances[22]) && (distances[9] < distances[23]) && (distances[9] < distances[24]) && (distances[9] < distances[25]) && (distances[9] < distances[26]) && (distances[9] < distances[27]) && (distances[9] < distances[28]) && (distances[9] < distances[29]) && (distances[9] < distances[30]) && (distances[9] < distances[31]) && (distances[9] < distances[32]) && (distances[9] < distances[33]) && (distances[9] < distances[34]) && (distances[9] < distances[35]) && (distances[9] < distances[36]) && (distances[9] < distances[37]) && (distances[9] < distances[38]) && (distances[9] < distances[39]) && (distances[9] < distances[40]) && (distances[9] < distances[41]) && (distances[9] < distances[42]) && (distances[9] < distances[43]) && (distances[9] < distances[44]) && (distances[9] < distances[45]) && (distances[9] < distances[46]) && (distances[9] < distances[47]) && (distances[9] < distances[48]) && (distances[9] < distances[49]) && (distances[9] < distances[50]) && (distances[9] < distances[51]) && (distances[9] < distances[52]) && (distances[9] < distances[53]) && (distances[9] < distances[54]) && (distances[9] < distances[55]) && (distances[9] < distances[56]) && (distances[9] < distances[57]) && (distances[9] < distances[58]) && (distances[9] < distances[59]) && (distances[9] < distances[60]) && (distances[9] < distances[61]) && (distances[9] < distances[62]) && (distances[9] < distances[63]) && (distances[9] < distances[64]) && (distances[9] < distances[65]) && (distances[9] < distances[66]) && (distances[9] < distances[67]) && (distances[9] < distances[68]) && (distances[9] < distances[69]) && (distances[9] < distances[70]) && (distances[9] < distances[71]) && (distances[9] < distances[72]) && (distances[9] < distances[73]) && (distances[9] < distances[74]) && (distances[9] < distances[75]) && (distances[9] < distances[76]) && (distances[9] < distances[77]) && (distances[9] < distances[78]) && (distances[9] < distances[79]) && (distances[9] < distances[80]) && (distances[9] < distances[81]) && (distances[9] < distances[82]) && (distances[9] < distances[83]) && (distances[9] < distances[84]) && (distances[9] < distances[85]) && (distances[9] < distances[86]) && (distances[9] < distances[87]) && (distances[9] < distances[88]) && (distances[9] < distances[89])) begin
        dout <= 9;
      end else if((distances[10] < distances[11]) && (distances[10] < distances[12]) && (distances[10] < distances[13]) && (distances[10] < distances[14]) && (distances[10] < distances[15]) && (distances[10] < distances[16]) && (distances[10] < distances[17]) && (distances[10] < distances[18]) && (distances[10] < distances[19]) && (distances[10] < distances[20]) && (distances[10] < distances[21]) && (distances[10] < distances[22]) && (distances[10] < distances[23]) && (distances[10] < distances[24]) && (distances[10] < distances[25]) && (distances[10] < distances[26]) && (distances[10] < distances[27]) && (distances[10] < distances[28]) && (distances[10] < distances[29]) && (distances[10] < distances[30]) && (distances[10] < distances[31]) && (distances[10] < distances[32]) && (distances[10] < distances[33]) && (distances[10] < distances[34]) && (distances[10] < distances[35]) && (distances[10] < distances[36]) && (distances[10] < distances[37]) && (distances[10] < distances[38]) && (distances[10] < distances[39]) && (distances[10] < distances[40]) && (distances[10] < distances[41]) && (distances[10] < distances[42]) && (distances[10] < distances[43]) && (distances[10] < distances[44]) && (distances[10] < distances[45]) && (distances[10] < distances[46]) && (distances[10] < distances[47]) && (distances[10] < distances[48]) && (distances[10] < distances[49]) && (distances[10] < distances[50]) && (distances[10] < distances[51]) && (distances[10] < distances[52]) && (distances[10] < distances[53]) && (distances[10] < distances[54]) && (distances[10] < distances[55]) && (distances[10] < distances[56]) && (distances[10] < distances[57]) && (distances[10] < distances[58]) && (distances[10] < distances[59]) && (distances[10] < distances[60]) && (distances[10] < distances[61]) && (distances[10] < distances[62]) && (distances[10] < distances[63]) && (distances[10] < distances[64]) && (distances[10] < distances[65]) && (distances[10] < distances[66]) && (distances[10] < distances[67]) && (distances[10] < distances[68]) && (distances[10] < distances[69]) && (distances[10] < distances[70]) && (distances[10] < distances[71]) && (distances[10] < distances[72]) && (distances[10] < distances[73]) && (distances[10] < distances[74]) && (distances[10] < distances[75]) && (distances[10] < distances[76]) && (distances[10] < distances[77]) && (distances[10] < distances[78]) && (distances[10] < distances[79]) && (distances[10] < distances[80]) && (distances[10] < distances[81]) && (distances[10] < distances[82]) && (distances[10] < distances[83]) && (distances[10] < distances[84]) && (distances[10] < distances[85]) && (distances[10] < distances[86]) && (distances[10] < distances[87]) && (distances[10] < distances[88]) && (distances[10] < distances[89])) begin
        dout <= 10;
      end else if((distances[11] < distances[12]) && (distances[11] < distances[13]) && (distances[11] < distances[14]) && (distances[11] < distances[15]) && (distances[11] < distances[16]) && (distances[11] < distances[17]) && (distances[11] < distances[18]) && (distances[11] < distances[19]) && (distances[11] < distances[20]) && (distances[11] < distances[21]) && (distances[11] < distances[22]) && (distances[11] < distances[23]) && (distances[11] < distances[24]) && (distances[11] < distances[25]) && (distances[11] < distances[26]) && (distances[11] < distances[27]) && (distances[11] < distances[28]) && (distances[11] < distances[29]) && (distances[11] < distances[30]) && (distances[11] < distances[31]) && (distances[11] < distances[32]) && (distances[11] < distances[33]) && (distances[11] < distances[34]) && (distances[11] < distances[35]) && (distances[11] < distances[36]) && (distances[11] < distances[37]) && (distances[11] < distances[38]) && (distances[11] < distances[39]) && (distances[11] < distances[40]) && (distances[11] < distances[41]) && (distances[11] < distances[42]) && (distances[11] < distances[43]) && (distances[11] < distances[44]) && (distances[11] < distances[45]) && (distances[11] < distances[46]) && (distances[11] < distances[47]) && (distances[11] < distances[48]) && (distances[11] < distances[49]) && (distances[11] < distances[50]) && (distances[11] < distances[51]) && (distances[11] < distances[52]) && (distances[11] < distances[53]) && (distances[11] < distances[54]) && (distances[11] < distances[55]) && (distances[11] < distances[56]) && (distances[11] < distances[57]) && (distances[11] < distances[58]) && (distances[11] < distances[59]) && (distances[11] < distances[60]) && (distances[11] < distances[61]) && (distances[11] < distances[62]) && (distances[11] < distances[63]) && (distances[11] < distances[64]) && (distances[11] < distances[65]) && (distances[11] < distances[66]) && (distances[11] < distances[67]) && (distances[11] < distances[68]) && (distances[11] < distances[69]) && (distances[11] < distances[70]) && (distances[11] < distances[71]) && (distances[11] < distances[72]) && (distances[11] < distances[73]) && (distances[11] < distances[74]) && (distances[11] < distances[75]) && (distances[11] < distances[76]) && (distances[11] < distances[77]) && (distances[11] < distances[78]) && (distances[11] < distances[79]) && (distances[11] < distances[80]) && (distances[11] < distances[81]) && (distances[11] < distances[82]) && (distances[11] < distances[83]) && (distances[11] < distances[84]) && (distances[11] < distances[85]) && (distances[11] < distances[86]) && (distances[11] < distances[87]) && (distances[11] < distances[88]) && (distances[11] < distances[89])) begin
        dout <= 11;
      end else if((distances[12] < distances[13]) && (distances[12] < distances[14]) && (distances[12] < distances[15]) && (distances[12] < distances[16]) && (distances[12] < distances[17]) && (distances[12] < distances[18]) && (distances[12] < distances[19]) && (distances[12] < distances[20]) && (distances[12] < distances[21]) && (distances[12] < distances[22]) && (distances[12] < distances[23]) && (distances[12] < distances[24]) && (distances[12] < distances[25]) && (distances[12] < distances[26]) && (distances[12] < distances[27]) && (distances[12] < distances[28]) && (distances[12] < distances[29]) && (distances[12] < distances[30]) && (distances[12] < distances[31]) && (distances[12] < distances[32]) && (distances[12] < distances[33]) && (distances[12] < distances[34]) && (distances[12] < distances[35]) && (distances[12] < distances[36]) && (distances[12] < distances[37]) && (distances[12] < distances[38]) && (distances[12] < distances[39]) && (distances[12] < distances[40]) && (distances[12] < distances[41]) && (distances[12] < distances[42]) && (distances[12] < distances[43]) && (distances[12] < distances[44]) && (distances[12] < distances[45]) && (distances[12] < distances[46]) && (distances[12] < distances[47]) && (distances[12] < distances[48]) && (distances[12] < distances[49]) && (distances[12] < distances[50]) && (distances[12] < distances[51]) && (distances[12] < distances[52]) && (distances[12] < distances[53]) && (distances[12] < distances[54]) && (distances[12] < distances[55]) && (distances[12] < distances[56]) && (distances[12] < distances[57]) && (distances[12] < distances[58]) && (distances[12] < distances[59]) && (distances[12] < distances[60]) && (distances[12] < distances[61]) && (distances[12] < distances[62]) && (distances[12] < distances[63]) && (distances[12] < distances[64]) && (distances[12] < distances[65]) && (distances[12] < distances[66]) && (distances[12] < distances[67]) && (distances[12] < distances[68]) && (distances[12] < distances[69]) && (distances[12] < distances[70]) && (distances[12] < distances[71]) && (distances[12] < distances[72]) && (distances[12] < distances[73]) && (distances[12] < distances[74]) && (distances[12] < distances[75]) && (distances[12] < distances[76]) && (distances[12] < distances[77]) && (distances[12] < distances[78]) && (distances[12] < distances[79]) && (distances[12] < distances[80]) && (distances[12] < distances[81]) && (distances[12] < distances[82]) && (distances[12] < distances[83]) && (distances[12] < distances[84]) && (distances[12] < distances[85]) && (distances[12] < distances[86]) && (distances[12] < distances[87]) && (distances[12] < distances[88]) && (distances[12] < distances[89])) begin
        dout <= 12;
      end else if((distances[13] < distances[14]) && (distances[13] < distances[15]) && (distances[13] < distances[16]) && (distances[13] < distances[17]) && (distances[13] < distances[18]) && (distances[13] < distances[19]) && (distances[13] < distances[20]) && (distances[13] < distances[21]) && (distances[13] < distances[22]) && (distances[13] < distances[23]) && (distances[13] < distances[24]) && (distances[13] < distances[25]) && (distances[13] < distances[26]) && (distances[13] < distances[27]) && (distances[13] < distances[28]) && (distances[13] < distances[29]) && (distances[13] < distances[30]) && (distances[13] < distances[31]) && (distances[13] < distances[32]) && (distances[13] < distances[33]) && (distances[13] < distances[34]) && (distances[13] < distances[35]) && (distances[13] < distances[36]) && (distances[13] < distances[37]) && (distances[13] < distances[38]) && (distances[13] < distances[39]) && (distances[13] < distances[40]) && (distances[13] < distances[41]) && (distances[13] < distances[42]) && (distances[13] < distances[43]) && (distances[13] < distances[44]) && (distances[13] < distances[45]) && (distances[13] < distances[46]) && (distances[13] < distances[47]) && (distances[13] < distances[48]) && (distances[13] < distances[49]) && (distances[13] < distances[50]) && (distances[13] < distances[51]) && (distances[13] < distances[52]) && (distances[13] < distances[53]) && (distances[13] < distances[54]) && (distances[13] < distances[55]) && (distances[13] < distances[56]) && (distances[13] < distances[57]) && (distances[13] < distances[58]) && (distances[13] < distances[59]) && (distances[13] < distances[60]) && (distances[13] < distances[61]) && (distances[13] < distances[62]) && (distances[13] < distances[63]) && (distances[13] < distances[64]) && (distances[13] < distances[65]) && (distances[13] < distances[66]) && (distances[13] < distances[67]) && (distances[13] < distances[68]) && (distances[13] < distances[69]) && (distances[13] < distances[70]) && (distances[13] < distances[71]) && (distances[13] < distances[72]) && (distances[13] < distances[73]) && (distances[13] < distances[74]) && (distances[13] < distances[75]) && (distances[13] < distances[76]) && (distances[13] < distances[77]) && (distances[13] < distances[78]) && (distances[13] < distances[79]) && (distances[13] < distances[80]) && (distances[13] < distances[81]) && (distances[13] < distances[82]) && (distances[13] < distances[83]) && (distances[13] < distances[84]) && (distances[13] < distances[85]) && (distances[13] < distances[86]) && (distances[13] < distances[87]) && (distances[13] < distances[88]) && (distances[13] < distances[89])) begin
        dout <= 13;
      end else if((distances[14] < distances[15]) && (distances[14] < distances[16]) && (distances[14] < distances[17]) && (distances[14] < distances[18]) && (distances[14] < distances[19]) && (distances[14] < distances[20]) && (distances[14] < distances[21]) && (distances[14] < distances[22]) && (distances[14] < distances[23]) && (distances[14] < distances[24]) && (distances[14] < distances[25]) && (distances[14] < distances[26]) && (distances[14] < distances[27]) && (distances[14] < distances[28]) && (distances[14] < distances[29]) && (distances[14] < distances[30]) && (distances[14] < distances[31]) && (distances[14] < distances[32]) && (distances[14] < distances[33]) && (distances[14] < distances[34]) && (distances[14] < distances[35]) && (distances[14] < distances[36]) && (distances[14] < distances[37]) && (distances[14] < distances[38]) && (distances[14] < distances[39]) && (distances[14] < distances[40]) && (distances[14] < distances[41]) && (distances[14] < distances[42]) && (distances[14] < distances[43]) && (distances[14] < distances[44]) && (distances[14] < distances[45]) && (distances[14] < distances[46]) && (distances[14] < distances[47]) && (distances[14] < distances[48]) && (distances[14] < distances[49]) && (distances[14] < distances[50]) && (distances[14] < distances[51]) && (distances[14] < distances[52]) && (distances[14] < distances[53]) && (distances[14] < distances[54]) && (distances[14] < distances[55]) && (distances[14] < distances[56]) && (distances[14] < distances[57]) && (distances[14] < distances[58]) && (distances[14] < distances[59]) && (distances[14] < distances[60]) && (distances[14] < distances[61]) && (distances[14] < distances[62]) && (distances[14] < distances[63]) && (distances[14] < distances[64]) && (distances[14] < distances[65]) && (distances[14] < distances[66]) && (distances[14] < distances[67]) && (distances[14] < distances[68]) && (distances[14] < distances[69]) && (distances[14] < distances[70]) && (distances[14] < distances[71]) && (distances[14] < distances[72]) && (distances[14] < distances[73]) && (distances[14] < distances[74]) && (distances[14] < distances[75]) && (distances[14] < distances[76]) && (distances[14] < distances[77]) && (distances[14] < distances[78]) && (distances[14] < distances[79]) && (distances[14] < distances[80]) && (distances[14] < distances[81]) && (distances[14] < distances[82]) && (distances[14] < distances[83]) && (distances[14] < distances[84]) && (distances[14] < distances[85]) && (distances[14] < distances[86]) && (distances[14] < distances[87]) && (distances[14] < distances[88]) && (distances[14] < distances[89])) begin
        dout <= 14;
      end else if((distances[15] < distances[16]) && (distances[15] < distances[17]) && (distances[15] < distances[18]) && (distances[15] < distances[19]) && (distances[15] < distances[20]) && (distances[15] < distances[21]) && (distances[15] < distances[22]) && (distances[15] < distances[23]) && (distances[15] < distances[24]) && (distances[15] < distances[25]) && (distances[15] < distances[26]) && (distances[15] < distances[27]) && (distances[15] < distances[28]) && (distances[15] < distances[29]) && (distances[15] < distances[30]) && (distances[15] < distances[31]) && (distances[15] < distances[32]) && (distances[15] < distances[33]) && (distances[15] < distances[34]) && (distances[15] < distances[35]) && (distances[15] < distances[36]) && (distances[15] < distances[37]) && (distances[15] < distances[38]) && (distances[15] < distances[39]) && (distances[15] < distances[40]) && (distances[15] < distances[41]) && (distances[15] < distances[42]) && (distances[15] < distances[43]) && (distances[15] < distances[44]) && (distances[15] < distances[45]) && (distances[15] < distances[46]) && (distances[15] < distances[47]) && (distances[15] < distances[48]) && (distances[15] < distances[49]) && (distances[15] < distances[50]) && (distances[15] < distances[51]) && (distances[15] < distances[52]) && (distances[15] < distances[53]) && (distances[15] < distances[54]) && (distances[15] < distances[55]) && (distances[15] < distances[56]) && (distances[15] < distances[57]) && (distances[15] < distances[58]) && (distances[15] < distances[59]) && (distances[15] < distances[60]) && (distances[15] < distances[61]) && (distances[15] < distances[62]) && (distances[15] < distances[63]) && (distances[15] < distances[64]) && (distances[15] < distances[65]) && (distances[15] < distances[66]) && (distances[15] < distances[67]) && (distances[15] < distances[68]) && (distances[15] < distances[69]) && (distances[15] < distances[70]) && (distances[15] < distances[71]) && (distances[15] < distances[72]) && (distances[15] < distances[73]) && (distances[15] < distances[74]) && (distances[15] < distances[75]) && (distances[15] < distances[76]) && (distances[15] < distances[77]) && (distances[15] < distances[78]) && (distances[15] < distances[79]) && (distances[15] < distances[80]) && (distances[15] < distances[81]) && (distances[15] < distances[82]) && (distances[15] < distances[83]) && (distances[15] < distances[84]) && (distances[15] < distances[85]) && (distances[15] < distances[86]) && (distances[15] < distances[87]) && (distances[15] < distances[88]) && (distances[15] < distances[89])) begin
        dout <= 15;
      end else if((distances[16] < distances[17]) && (distances[16] < distances[18]) && (distances[16] < distances[19]) && (distances[16] < distances[20]) && (distances[16] < distances[21]) && (distances[16] < distances[22]) && (distances[16] < distances[23]) && (distances[16] < distances[24]) && (distances[16] < distances[25]) && (distances[16] < distances[26]) && (distances[16] < distances[27]) && (distances[16] < distances[28]) && (distances[16] < distances[29]) && (distances[16] < distances[30]) && (distances[16] < distances[31]) && (distances[16] < distances[32]) && (distances[16] < distances[33]) && (distances[16] < distances[34]) && (distances[16] < distances[35]) && (distances[16] < distances[36]) && (distances[16] < distances[37]) && (distances[16] < distances[38]) && (distances[16] < distances[39]) && (distances[16] < distances[40]) && (distances[16] < distances[41]) && (distances[16] < distances[42]) && (distances[16] < distances[43]) && (distances[16] < distances[44]) && (distances[16] < distances[45]) && (distances[16] < distances[46]) && (distances[16] < distances[47]) && (distances[16] < distances[48]) && (distances[16] < distances[49]) && (distances[16] < distances[50]) && (distances[16] < distances[51]) && (distances[16] < distances[52]) && (distances[16] < distances[53]) && (distances[16] < distances[54]) && (distances[16] < distances[55]) && (distances[16] < distances[56]) && (distances[16] < distances[57]) && (distances[16] < distances[58]) && (distances[16] < distances[59]) && (distances[16] < distances[60]) && (distances[16] < distances[61]) && (distances[16] < distances[62]) && (distances[16] < distances[63]) && (distances[16] < distances[64]) && (distances[16] < distances[65]) && (distances[16] < distances[66]) && (distances[16] < distances[67]) && (distances[16] < distances[68]) && (distances[16] < distances[69]) && (distances[16] < distances[70]) && (distances[16] < distances[71]) && (distances[16] < distances[72]) && (distances[16] < distances[73]) && (distances[16] < distances[74]) && (distances[16] < distances[75]) && (distances[16] < distances[76]) && (distances[16] < distances[77]) && (distances[16] < distances[78]) && (distances[16] < distances[79]) && (distances[16] < distances[80]) && (distances[16] < distances[81]) && (distances[16] < distances[82]) && (distances[16] < distances[83]) && (distances[16] < distances[84]) && (distances[16] < distances[85]) && (distances[16] < distances[86]) && (distances[16] < distances[87]) && (distances[16] < distances[88]) && (distances[16] < distances[89])) begin
        dout <= 16;
      end else if((distances[17] < distances[18]) && (distances[17] < distances[19]) && (distances[17] < distances[20]) && (distances[17] < distances[21]) && (distances[17] < distances[22]) && (distances[17] < distances[23]) && (distances[17] < distances[24]) && (distances[17] < distances[25]) && (distances[17] < distances[26]) && (distances[17] < distances[27]) && (distances[17] < distances[28]) && (distances[17] < distances[29]) && (distances[17] < distances[30]) && (distances[17] < distances[31]) && (distances[17] < distances[32]) && (distances[17] < distances[33]) && (distances[17] < distances[34]) && (distances[17] < distances[35]) && (distances[17] < distances[36]) && (distances[17] < distances[37]) && (distances[17] < distances[38]) && (distances[17] < distances[39]) && (distances[17] < distances[40]) && (distances[17] < distances[41]) && (distances[17] < distances[42]) && (distances[17] < distances[43]) && (distances[17] < distances[44]) && (distances[17] < distances[45]) && (distances[17] < distances[46]) && (distances[17] < distances[47]) && (distances[17] < distances[48]) && (distances[17] < distances[49]) && (distances[17] < distances[50]) && (distances[17] < distances[51]) && (distances[17] < distances[52]) && (distances[17] < distances[53]) && (distances[17] < distances[54]) && (distances[17] < distances[55]) && (distances[17] < distances[56]) && (distances[17] < distances[57]) && (distances[17] < distances[58]) && (distances[17] < distances[59]) && (distances[17] < distances[60]) && (distances[17] < distances[61]) && (distances[17] < distances[62]) && (distances[17] < distances[63]) && (distances[17] < distances[64]) && (distances[17] < distances[65]) && (distances[17] < distances[66]) && (distances[17] < distances[67]) && (distances[17] < distances[68]) && (distances[17] < distances[69]) && (distances[17] < distances[70]) && (distances[17] < distances[71]) && (distances[17] < distances[72]) && (distances[17] < distances[73]) && (distances[17] < distances[74]) && (distances[17] < distances[75]) && (distances[17] < distances[76]) && (distances[17] < distances[77]) && (distances[17] < distances[78]) && (distances[17] < distances[79]) && (distances[17] < distances[80]) && (distances[17] < distances[81]) && (distances[17] < distances[82]) && (distances[17] < distances[83]) && (distances[17] < distances[84]) && (distances[17] < distances[85]) && (distances[17] < distances[86]) && (distances[17] < distances[87]) && (distances[17] < distances[88]) && (distances[17] < distances[89])) begin
        dout <= 17;
      end else if((distances[18] < distances[19]) && (distances[18] < distances[20]) && (distances[18] < distances[21]) && (distances[18] < distances[22]) && (distances[18] < distances[23]) && (distances[18] < distances[24]) && (distances[18] < distances[25]) && (distances[18] < distances[26]) && (distances[18] < distances[27]) && (distances[18] < distances[28]) && (distances[18] < distances[29]) && (distances[18] < distances[30]) && (distances[18] < distances[31]) && (distances[18] < distances[32]) && (distances[18] < distances[33]) && (distances[18] < distances[34]) && (distances[18] < distances[35]) && (distances[18] < distances[36]) && (distances[18] < distances[37]) && (distances[18] < distances[38]) && (distances[18] < distances[39]) && (distances[18] < distances[40]) && (distances[18] < distances[41]) && (distances[18] < distances[42]) && (distances[18] < distances[43]) && (distances[18] < distances[44]) && (distances[18] < distances[45]) && (distances[18] < distances[46]) && (distances[18] < distances[47]) && (distances[18] < distances[48]) && (distances[18] < distances[49]) && (distances[18] < distances[50]) && (distances[18] < distances[51]) && (distances[18] < distances[52]) && (distances[18] < distances[53]) && (distances[18] < distances[54]) && (distances[18] < distances[55]) && (distances[18] < distances[56]) && (distances[18] < distances[57]) && (distances[18] < distances[58]) && (distances[18] < distances[59]) && (distances[18] < distances[60]) && (distances[18] < distances[61]) && (distances[18] < distances[62]) && (distances[18] < distances[63]) && (distances[18] < distances[64]) && (distances[18] < distances[65]) && (distances[18] < distances[66]) && (distances[18] < distances[67]) && (distances[18] < distances[68]) && (distances[18] < distances[69]) && (distances[18] < distances[70]) && (distances[18] < distances[71]) && (distances[18] < distances[72]) && (distances[18] < distances[73]) && (distances[18] < distances[74]) && (distances[18] < distances[75]) && (distances[18] < distances[76]) && (distances[18] < distances[77]) && (distances[18] < distances[78]) && (distances[18] < distances[79]) && (distances[18] < distances[80]) && (distances[18] < distances[81]) && (distances[18] < distances[82]) && (distances[18] < distances[83]) && (distances[18] < distances[84]) && (distances[18] < distances[85]) && (distances[18] < distances[86]) && (distances[18] < distances[87]) && (distances[18] < distances[88]) && (distances[18] < distances[89])) begin
        dout <= 18;
      end else if((distances[19] < distances[20]) && (distances[19] < distances[21]) && (distances[19] < distances[22]) && (distances[19] < distances[23]) && (distances[19] < distances[24]) && (distances[19] < distances[25]) && (distances[19] < distances[26]) && (distances[19] < distances[27]) && (distances[19] < distances[28]) && (distances[19] < distances[29]) && (distances[19] < distances[30]) && (distances[19] < distances[31]) && (distances[19] < distances[32]) && (distances[19] < distances[33]) && (distances[19] < distances[34]) && (distances[19] < distances[35]) && (distances[19] < distances[36]) && (distances[19] < distances[37]) && (distances[19] < distances[38]) && (distances[19] < distances[39]) && (distances[19] < distances[40]) && (distances[19] < distances[41]) && (distances[19] < distances[42]) && (distances[19] < distances[43]) && (distances[19] < distances[44]) && (distances[19] < distances[45]) && (distances[19] < distances[46]) && (distances[19] < distances[47]) && (distances[19] < distances[48]) && (distances[19] < distances[49]) && (distances[19] < distances[50]) && (distances[19] < distances[51]) && (distances[19] < distances[52]) && (distances[19] < distances[53]) && (distances[19] < distances[54]) && (distances[19] < distances[55]) && (distances[19] < distances[56]) && (distances[19] < distances[57]) && (distances[19] < distances[58]) && (distances[19] < distances[59]) && (distances[19] < distances[60]) && (distances[19] < distances[61]) && (distances[19] < distances[62]) && (distances[19] < distances[63]) && (distances[19] < distances[64]) && (distances[19] < distances[65]) && (distances[19] < distances[66]) && (distances[19] < distances[67]) && (distances[19] < distances[68]) && (distances[19] < distances[69]) && (distances[19] < distances[70]) && (distances[19] < distances[71]) && (distances[19] < distances[72]) && (distances[19] < distances[73]) && (distances[19] < distances[74]) && (distances[19] < distances[75]) && (distances[19] < distances[76]) && (distances[19] < distances[77]) && (distances[19] < distances[78]) && (distances[19] < distances[79]) && (distances[19] < distances[80]) && (distances[19] < distances[81]) && (distances[19] < distances[82]) && (distances[19] < distances[83]) && (distances[19] < distances[84]) && (distances[19] < distances[85]) && (distances[19] < distances[86]) && (distances[19] < distances[87]) && (distances[19] < distances[88]) && (distances[19] < distances[89])) begin
        dout <= 19;
      end else if((distances[20] < distances[21]) && (distances[20] < distances[22]) && (distances[20] < distances[23]) && (distances[20] < distances[24]) && (distances[20] < distances[25]) && (distances[20] < distances[26]) && (distances[20] < distances[27]) && (distances[20] < distances[28]) && (distances[20] < distances[29]) && (distances[20] < distances[30]) && (distances[20] < distances[31]) && (distances[20] < distances[32]) && (distances[20] < distances[33]) && (distances[20] < distances[34]) && (distances[20] < distances[35]) && (distances[20] < distances[36]) && (distances[20] < distances[37]) && (distances[20] < distances[38]) && (distances[20] < distances[39]) && (distances[20] < distances[40]) && (distances[20] < distances[41]) && (distances[20] < distances[42]) && (distances[20] < distances[43]) && (distances[20] < distances[44]) && (distances[20] < distances[45]) && (distances[20] < distances[46]) && (distances[20] < distances[47]) && (distances[20] < distances[48]) && (distances[20] < distances[49]) && (distances[20] < distances[50]) && (distances[20] < distances[51]) && (distances[20] < distances[52]) && (distances[20] < distances[53]) && (distances[20] < distances[54]) && (distances[20] < distances[55]) && (distances[20] < distances[56]) && (distances[20] < distances[57]) && (distances[20] < distances[58]) && (distances[20] < distances[59]) && (distances[20] < distances[60]) && (distances[20] < distances[61]) && (distances[20] < distances[62]) && (distances[20] < distances[63]) && (distances[20] < distances[64]) && (distances[20] < distances[65]) && (distances[20] < distances[66]) && (distances[20] < distances[67]) && (distances[20] < distances[68]) && (distances[20] < distances[69]) && (distances[20] < distances[70]) && (distances[20] < distances[71]) && (distances[20] < distances[72]) && (distances[20] < distances[73]) && (distances[20] < distances[74]) && (distances[20] < distances[75]) && (distances[20] < distances[76]) && (distances[20] < distances[77]) && (distances[20] < distances[78]) && (distances[20] < distances[79]) && (distances[20] < distances[80]) && (distances[20] < distances[81]) && (distances[20] < distances[82]) && (distances[20] < distances[83]) && (distances[20] < distances[84]) && (distances[20] < distances[85]) && (distances[20] < distances[86]) && (distances[20] < distances[87]) && (distances[20] < distances[88]) && (distances[20] < distances[89])) begin
        dout <= 20;
      end else if((distances[21] < distances[22]) && (distances[21] < distances[23]) && (distances[21] < distances[24]) && (distances[21] < distances[25]) && (distances[21] < distances[26]) && (distances[21] < distances[27]) && (distances[21] < distances[28]) && (distances[21] < distances[29]) && (distances[21] < distances[30]) && (distances[21] < distances[31]) && (distances[21] < distances[32]) && (distances[21] < distances[33]) && (distances[21] < distances[34]) && (distances[21] < distances[35]) && (distances[21] < distances[36]) && (distances[21] < distances[37]) && (distances[21] < distances[38]) && (distances[21] < distances[39]) && (distances[21] < distances[40]) && (distances[21] < distances[41]) && (distances[21] < distances[42]) && (distances[21] < distances[43]) && (distances[21] < distances[44]) && (distances[21] < distances[45]) && (distances[21] < distances[46]) && (distances[21] < distances[47]) && (distances[21] < distances[48]) && (distances[21] < distances[49]) && (distances[21] < distances[50]) && (distances[21] < distances[51]) && (distances[21] < distances[52]) && (distances[21] < distances[53]) && (distances[21] < distances[54]) && (distances[21] < distances[55]) && (distances[21] < distances[56]) && (distances[21] < distances[57]) && (distances[21] < distances[58]) && (distances[21] < distances[59]) && (distances[21] < distances[60]) && (distances[21] < distances[61]) && (distances[21] < distances[62]) && (distances[21] < distances[63]) && (distances[21] < distances[64]) && (distances[21] < distances[65]) && (distances[21] < distances[66]) && (distances[21] < distances[67]) && (distances[21] < distances[68]) && (distances[21] < distances[69]) && (distances[21] < distances[70]) && (distances[21] < distances[71]) && (distances[21] < distances[72]) && (distances[21] < distances[73]) && (distances[21] < distances[74]) && (distances[21] < distances[75]) && (distances[21] < distances[76]) && (distances[21] < distances[77]) && (distances[21] < distances[78]) && (distances[21] < distances[79]) && (distances[21] < distances[80]) && (distances[21] < distances[81]) && (distances[21] < distances[82]) && (distances[21] < distances[83]) && (distances[21] < distances[84]) && (distances[21] < distances[85]) && (distances[21] < distances[86]) && (distances[21] < distances[87]) && (distances[21] < distances[88]) && (distances[21] < distances[89])) begin
        dout <= 21;
      end else if((distances[22] < distances[23]) && (distances[22] < distances[24]) && (distances[22] < distances[25]) && (distances[22] < distances[26]) && (distances[22] < distances[27]) && (distances[22] < distances[28]) && (distances[22] < distances[29]) && (distances[22] < distances[30]) && (distances[22] < distances[31]) && (distances[22] < distances[32]) && (distances[22] < distances[33]) && (distances[22] < distances[34]) && (distances[22] < distances[35]) && (distances[22] < distances[36]) && (distances[22] < distances[37]) && (distances[22] < distances[38]) && (distances[22] < distances[39]) && (distances[22] < distances[40]) && (distances[22] < distances[41]) && (distances[22] < distances[42]) && (distances[22] < distances[43]) && (distances[22] < distances[44]) && (distances[22] < distances[45]) && (distances[22] < distances[46]) && (distances[22] < distances[47]) && (distances[22] < distances[48]) && (distances[22] < distances[49]) && (distances[22] < distances[50]) && (distances[22] < distances[51]) && (distances[22] < distances[52]) && (distances[22] < distances[53]) && (distances[22] < distances[54]) && (distances[22] < distances[55]) && (distances[22] < distances[56]) && (distances[22] < distances[57]) && (distances[22] < distances[58]) && (distances[22] < distances[59]) && (distances[22] < distances[60]) && (distances[22] < distances[61]) && (distances[22] < distances[62]) && (distances[22] < distances[63]) && (distances[22] < distances[64]) && (distances[22] < distances[65]) && (distances[22] < distances[66]) && (distances[22] < distances[67]) && (distances[22] < distances[68]) && (distances[22] < distances[69]) && (distances[22] < distances[70]) && (distances[22] < distances[71]) && (distances[22] < distances[72]) && (distances[22] < distances[73]) && (distances[22] < distances[74]) && (distances[22] < distances[75]) && (distances[22] < distances[76]) && (distances[22] < distances[77]) && (distances[22] < distances[78]) && (distances[22] < distances[79]) && (distances[22] < distances[80]) && (distances[22] < distances[81]) && (distances[22] < distances[82]) && (distances[22] < distances[83]) && (distances[22] < distances[84]) && (distances[22] < distances[85]) && (distances[22] < distances[86]) && (distances[22] < distances[87]) && (distances[22] < distances[88]) && (distances[22] < distances[89])) begin
        dout <= 22;
      end else if((distances[23] < distances[24]) && (distances[23] < distances[25]) && (distances[23] < distances[26]) && (distances[23] < distances[27]) && (distances[23] < distances[28]) && (distances[23] < distances[29]) && (distances[23] < distances[30]) && (distances[23] < distances[31]) && (distances[23] < distances[32]) && (distances[23] < distances[33]) && (distances[23] < distances[34]) && (distances[23] < distances[35]) && (distances[23] < distances[36]) && (distances[23] < distances[37]) && (distances[23] < distances[38]) && (distances[23] < distances[39]) && (distances[23] < distances[40]) && (distances[23] < distances[41]) && (distances[23] < distances[42]) && (distances[23] < distances[43]) && (distances[23] < distances[44]) && (distances[23] < distances[45]) && (distances[23] < distances[46]) && (distances[23] < distances[47]) && (distances[23] < distances[48]) && (distances[23] < distances[49]) && (distances[23] < distances[50]) && (distances[23] < distances[51]) && (distances[23] < distances[52]) && (distances[23] < distances[53]) && (distances[23] < distances[54]) && (distances[23] < distances[55]) && (distances[23] < distances[56]) && (distances[23] < distances[57]) && (distances[23] < distances[58]) && (distances[23] < distances[59]) && (distances[23] < distances[60]) && (distances[23] < distances[61]) && (distances[23] < distances[62]) && (distances[23] < distances[63]) && (distances[23] < distances[64]) && (distances[23] < distances[65]) && (distances[23] < distances[66]) && (distances[23] < distances[67]) && (distances[23] < distances[68]) && (distances[23] < distances[69]) && (distances[23] < distances[70]) && (distances[23] < distances[71]) && (distances[23] < distances[72]) && (distances[23] < distances[73]) && (distances[23] < distances[74]) && (distances[23] < distances[75]) && (distances[23] < distances[76]) && (distances[23] < distances[77]) && (distances[23] < distances[78]) && (distances[23] < distances[79]) && (distances[23] < distances[80]) && (distances[23] < distances[81]) && (distances[23] < distances[82]) && (distances[23] < distances[83]) && (distances[23] < distances[84]) && (distances[23] < distances[85]) && (distances[23] < distances[86]) && (distances[23] < distances[87]) && (distances[23] < distances[88]) && (distances[23] < distances[89])) begin
        dout <= 23;
      end else if((distances[24] < distances[25]) && (distances[24] < distances[26]) && (distances[24] < distances[27]) && (distances[24] < distances[28]) && (distances[24] < distances[29]) && (distances[24] < distances[30]) && (distances[24] < distances[31]) && (distances[24] < distances[32]) && (distances[24] < distances[33]) && (distances[24] < distances[34]) && (distances[24] < distances[35]) && (distances[24] < distances[36]) && (distances[24] < distances[37]) && (distances[24] < distances[38]) && (distances[24] < distances[39]) && (distances[24] < distances[40]) && (distances[24] < distances[41]) && (distances[24] < distances[42]) && (distances[24] < distances[43]) && (distances[24] < distances[44]) && (distances[24] < distances[45]) && (distances[24] < distances[46]) && (distances[24] < distances[47]) && (distances[24] < distances[48]) && (distances[24] < distances[49]) && (distances[24] < distances[50]) && (distances[24] < distances[51]) && (distances[24] < distances[52]) && (distances[24] < distances[53]) && (distances[24] < distances[54]) && (distances[24] < distances[55]) && (distances[24] < distances[56]) && (distances[24] < distances[57]) && (distances[24] < distances[58]) && (distances[24] < distances[59]) && (distances[24] < distances[60]) && (distances[24] < distances[61]) && (distances[24] < distances[62]) && (distances[24] < distances[63]) && (distances[24] < distances[64]) && (distances[24] < distances[65]) && (distances[24] < distances[66]) && (distances[24] < distances[67]) && (distances[24] < distances[68]) && (distances[24] < distances[69]) && (distances[24] < distances[70]) && (distances[24] < distances[71]) && (distances[24] < distances[72]) && (distances[24] < distances[73]) && (distances[24] < distances[74]) && (distances[24] < distances[75]) && (distances[24] < distances[76]) && (distances[24] < distances[77]) && (distances[24] < distances[78]) && (distances[24] < distances[79]) && (distances[24] < distances[80]) && (distances[24] < distances[81]) && (distances[24] < distances[82]) && (distances[24] < distances[83]) && (distances[24] < distances[84]) && (distances[24] < distances[85]) && (distances[24] < distances[86]) && (distances[24] < distances[87]) && (distances[24] < distances[88]) && (distances[24] < distances[89])) begin
        dout <= 24;
      end else if((distances[25] < distances[26]) && (distances[25] < distances[27]) && (distances[25] < distances[28]) && (distances[25] < distances[29]) && (distances[25] < distances[30]) && (distances[25] < distances[31]) && (distances[25] < distances[32]) && (distances[25] < distances[33]) && (distances[25] < distances[34]) && (distances[25] < distances[35]) && (distances[25] < distances[36]) && (distances[25] < distances[37]) && (distances[25] < distances[38]) && (distances[25] < distances[39]) && (distances[25] < distances[40]) && (distances[25] < distances[41]) && (distances[25] < distances[42]) && (distances[25] < distances[43]) && (distances[25] < distances[44]) && (distances[25] < distances[45]) && (distances[25] < distances[46]) && (distances[25] < distances[47]) && (distances[25] < distances[48]) && (distances[25] < distances[49]) && (distances[25] < distances[50]) && (distances[25] < distances[51]) && (distances[25] < distances[52]) && (distances[25] < distances[53]) && (distances[25] < distances[54]) && (distances[25] < distances[55]) && (distances[25] < distances[56]) && (distances[25] < distances[57]) && (distances[25] < distances[58]) && (distances[25] < distances[59]) && (distances[25] < distances[60]) && (distances[25] < distances[61]) && (distances[25] < distances[62]) && (distances[25] < distances[63]) && (distances[25] < distances[64]) && (distances[25] < distances[65]) && (distances[25] < distances[66]) && (distances[25] < distances[67]) && (distances[25] < distances[68]) && (distances[25] < distances[69]) && (distances[25] < distances[70]) && (distances[25] < distances[71]) && (distances[25] < distances[72]) && (distances[25] < distances[73]) && (distances[25] < distances[74]) && (distances[25] < distances[75]) && (distances[25] < distances[76]) && (distances[25] < distances[77]) && (distances[25] < distances[78]) && (distances[25] < distances[79]) && (distances[25] < distances[80]) && (distances[25] < distances[81]) && (distances[25] < distances[82]) && (distances[25] < distances[83]) && (distances[25] < distances[84]) && (distances[25] < distances[85]) && (distances[25] < distances[86]) && (distances[25] < distances[87]) && (distances[25] < distances[88]) && (distances[25] < distances[89])) begin
        dout <= 25;
      end else if((distances[26] < distances[27]) && (distances[26] < distances[28]) && (distances[26] < distances[29]) && (distances[26] < distances[30]) && (distances[26] < distances[31]) && (distances[26] < distances[32]) && (distances[26] < distances[33]) && (distances[26] < distances[34]) && (distances[26] < distances[35]) && (distances[26] < distances[36]) && (distances[26] < distances[37]) && (distances[26] < distances[38]) && (distances[26] < distances[39]) && (distances[26] < distances[40]) && (distances[26] < distances[41]) && (distances[26] < distances[42]) && (distances[26] < distances[43]) && (distances[26] < distances[44]) && (distances[26] < distances[45]) && (distances[26] < distances[46]) && (distances[26] < distances[47]) && (distances[26] < distances[48]) && (distances[26] < distances[49]) && (distances[26] < distances[50]) && (distances[26] < distances[51]) && (distances[26] < distances[52]) && (distances[26] < distances[53]) && (distances[26] < distances[54]) && (distances[26] < distances[55]) && (distances[26] < distances[56]) && (distances[26] < distances[57]) && (distances[26] < distances[58]) && (distances[26] < distances[59]) && (distances[26] < distances[60]) && (distances[26] < distances[61]) && (distances[26] < distances[62]) && (distances[26] < distances[63]) && (distances[26] < distances[64]) && (distances[26] < distances[65]) && (distances[26] < distances[66]) && (distances[26] < distances[67]) && (distances[26] < distances[68]) && (distances[26] < distances[69]) && (distances[26] < distances[70]) && (distances[26] < distances[71]) && (distances[26] < distances[72]) && (distances[26] < distances[73]) && (distances[26] < distances[74]) && (distances[26] < distances[75]) && (distances[26] < distances[76]) && (distances[26] < distances[77]) && (distances[26] < distances[78]) && (distances[26] < distances[79]) && (distances[26] < distances[80]) && (distances[26] < distances[81]) && (distances[26] < distances[82]) && (distances[26] < distances[83]) && (distances[26] < distances[84]) && (distances[26] < distances[85]) && (distances[26] < distances[86]) && (distances[26] < distances[87]) && (distances[26] < distances[88]) && (distances[26] < distances[89])) begin
        dout <= 26;
      end else if((distances[27] < distances[28]) && (distances[27] < distances[29]) && (distances[27] < distances[30]) && (distances[27] < distances[31]) && (distances[27] < distances[32]) && (distances[27] < distances[33]) && (distances[27] < distances[34]) && (distances[27] < distances[35]) && (distances[27] < distances[36]) && (distances[27] < distances[37]) && (distances[27] < distances[38]) && (distances[27] < distances[39]) && (distances[27] < distances[40]) && (distances[27] < distances[41]) && (distances[27] < distances[42]) && (distances[27] < distances[43]) && (distances[27] < distances[44]) && (distances[27] < distances[45]) && (distances[27] < distances[46]) && (distances[27] < distances[47]) && (distances[27] < distances[48]) && (distances[27] < distances[49]) && (distances[27] < distances[50]) && (distances[27] < distances[51]) && (distances[27] < distances[52]) && (distances[27] < distances[53]) && (distances[27] < distances[54]) && (distances[27] < distances[55]) && (distances[27] < distances[56]) && (distances[27] < distances[57]) && (distances[27] < distances[58]) && (distances[27] < distances[59]) && (distances[27] < distances[60]) && (distances[27] < distances[61]) && (distances[27] < distances[62]) && (distances[27] < distances[63]) && (distances[27] < distances[64]) && (distances[27] < distances[65]) && (distances[27] < distances[66]) && (distances[27] < distances[67]) && (distances[27] < distances[68]) && (distances[27] < distances[69]) && (distances[27] < distances[70]) && (distances[27] < distances[71]) && (distances[27] < distances[72]) && (distances[27] < distances[73]) && (distances[27] < distances[74]) && (distances[27] < distances[75]) && (distances[27] < distances[76]) && (distances[27] < distances[77]) && (distances[27] < distances[78]) && (distances[27] < distances[79]) && (distances[27] < distances[80]) && (distances[27] < distances[81]) && (distances[27] < distances[82]) && (distances[27] < distances[83]) && (distances[27] < distances[84]) && (distances[27] < distances[85]) && (distances[27] < distances[86]) && (distances[27] < distances[87]) && (distances[27] < distances[88]) && (distances[27] < distances[89])) begin
        dout <= 27;
      end else if((distances[28] < distances[29]) && (distances[28] < distances[30]) && (distances[28] < distances[31]) && (distances[28] < distances[32]) && (distances[28] < distances[33]) && (distances[28] < distances[34]) && (distances[28] < distances[35]) && (distances[28] < distances[36]) && (distances[28] < distances[37]) && (distances[28] < distances[38]) && (distances[28] < distances[39]) && (distances[28] < distances[40]) && (distances[28] < distances[41]) && (distances[28] < distances[42]) && (distances[28] < distances[43]) && (distances[28] < distances[44]) && (distances[28] < distances[45]) && (distances[28] < distances[46]) && (distances[28] < distances[47]) && (distances[28] < distances[48]) && (distances[28] < distances[49]) && (distances[28] < distances[50]) && (distances[28] < distances[51]) && (distances[28] < distances[52]) && (distances[28] < distances[53]) && (distances[28] < distances[54]) && (distances[28] < distances[55]) && (distances[28] < distances[56]) && (distances[28] < distances[57]) && (distances[28] < distances[58]) && (distances[28] < distances[59]) && (distances[28] < distances[60]) && (distances[28] < distances[61]) && (distances[28] < distances[62]) && (distances[28] < distances[63]) && (distances[28] < distances[64]) && (distances[28] < distances[65]) && (distances[28] < distances[66]) && (distances[28] < distances[67]) && (distances[28] < distances[68]) && (distances[28] < distances[69]) && (distances[28] < distances[70]) && (distances[28] < distances[71]) && (distances[28] < distances[72]) && (distances[28] < distances[73]) && (distances[28] < distances[74]) && (distances[28] < distances[75]) && (distances[28] < distances[76]) && (distances[28] < distances[77]) && (distances[28] < distances[78]) && (distances[28] < distances[79]) && (distances[28] < distances[80]) && (distances[28] < distances[81]) && (distances[28] < distances[82]) && (distances[28] < distances[83]) && (distances[28] < distances[84]) && (distances[28] < distances[85]) && (distances[28] < distances[86]) && (distances[28] < distances[87]) && (distances[28] < distances[88]) && (distances[28] < distances[89])) begin
        dout <= 28;
      end else if((distances[29] < distances[30]) && (distances[29] < distances[31]) && (distances[29] < distances[32]) && (distances[29] < distances[33]) && (distances[29] < distances[34]) && (distances[29] < distances[35]) && (distances[29] < distances[36]) && (distances[29] < distances[37]) && (distances[29] < distances[38]) && (distances[29] < distances[39]) && (distances[29] < distances[40]) && (distances[29] < distances[41]) && (distances[29] < distances[42]) && (distances[29] < distances[43]) && (distances[29] < distances[44]) && (distances[29] < distances[45]) && (distances[29] < distances[46]) && (distances[29] < distances[47]) && (distances[29] < distances[48]) && (distances[29] < distances[49]) && (distances[29] < distances[50]) && (distances[29] < distances[51]) && (distances[29] < distances[52]) && (distances[29] < distances[53]) && (distances[29] < distances[54]) && (distances[29] < distances[55]) && (distances[29] < distances[56]) && (distances[29] < distances[57]) && (distances[29] < distances[58]) && (distances[29] < distances[59]) && (distances[29] < distances[60]) && (distances[29] < distances[61]) && (distances[29] < distances[62]) && (distances[29] < distances[63]) && (distances[29] < distances[64]) && (distances[29] < distances[65]) && (distances[29] < distances[66]) && (distances[29] < distances[67]) && (distances[29] < distances[68]) && (distances[29] < distances[69]) && (distances[29] < distances[70]) && (distances[29] < distances[71]) && (distances[29] < distances[72]) && (distances[29] < distances[73]) && (distances[29] < distances[74]) && (distances[29] < distances[75]) && (distances[29] < distances[76]) && (distances[29] < distances[77]) && (distances[29] < distances[78]) && (distances[29] < distances[79]) && (distances[29] < distances[80]) && (distances[29] < distances[81]) && (distances[29] < distances[82]) && (distances[29] < distances[83]) && (distances[29] < distances[84]) && (distances[29] < distances[85]) && (distances[29] < distances[86]) && (distances[29] < distances[87]) && (distances[29] < distances[88]) && (distances[29] < distances[89])) begin
        dout <= 29;
      end else if((distances[30] < distances[31]) && (distances[30] < distances[32]) && (distances[30] < distances[33]) && (distances[30] < distances[34]) && (distances[30] < distances[35]) && (distances[30] < distances[36]) && (distances[30] < distances[37]) && (distances[30] < distances[38]) && (distances[30] < distances[39]) && (distances[30] < distances[40]) && (distances[30] < distances[41]) && (distances[30] < distances[42]) && (distances[30] < distances[43]) && (distances[30] < distances[44]) && (distances[30] < distances[45]) && (distances[30] < distances[46]) && (distances[30] < distances[47]) && (distances[30] < distances[48]) && (distances[30] < distances[49]) && (distances[30] < distances[50]) && (distances[30] < distances[51]) && (distances[30] < distances[52]) && (distances[30] < distances[53]) && (distances[30] < distances[54]) && (distances[30] < distances[55]) && (distances[30] < distances[56]) && (distances[30] < distances[57]) && (distances[30] < distances[58]) && (distances[30] < distances[59]) && (distances[30] < distances[60]) && (distances[30] < distances[61]) && (distances[30] < distances[62]) && (distances[30] < distances[63]) && (distances[30] < distances[64]) && (distances[30] < distances[65]) && (distances[30] < distances[66]) && (distances[30] < distances[67]) && (distances[30] < distances[68]) && (distances[30] < distances[69]) && (distances[30] < distances[70]) && (distances[30] < distances[71]) && (distances[30] < distances[72]) && (distances[30] < distances[73]) && (distances[30] < distances[74]) && (distances[30] < distances[75]) && (distances[30] < distances[76]) && (distances[30] < distances[77]) && (distances[30] < distances[78]) && (distances[30] < distances[79]) && (distances[30] < distances[80]) && (distances[30] < distances[81]) && (distances[30] < distances[82]) && (distances[30] < distances[83]) && (distances[30] < distances[84]) && (distances[30] < distances[85]) && (distances[30] < distances[86]) && (distances[30] < distances[87]) && (distances[30] < distances[88]) && (distances[30] < distances[89])) begin
        dout <= 30;
      end else if((distances[31] < distances[32]) && (distances[31] < distances[33]) && (distances[31] < distances[34]) && (distances[31] < distances[35]) && (distances[31] < distances[36]) && (distances[31] < distances[37]) && (distances[31] < distances[38]) && (distances[31] < distances[39]) && (distances[31] < distances[40]) && (distances[31] < distances[41]) && (distances[31] < distances[42]) && (distances[31] < distances[43]) && (distances[31] < distances[44]) && (distances[31] < distances[45]) && (distances[31] < distances[46]) && (distances[31] < distances[47]) && (distances[31] < distances[48]) && (distances[31] < distances[49]) && (distances[31] < distances[50]) && (distances[31] < distances[51]) && (distances[31] < distances[52]) && (distances[31] < distances[53]) && (distances[31] < distances[54]) && (distances[31] < distances[55]) && (distances[31] < distances[56]) && (distances[31] < distances[57]) && (distances[31] < distances[58]) && (distances[31] < distances[59]) && (distances[31] < distances[60]) && (distances[31] < distances[61]) && (distances[31] < distances[62]) && (distances[31] < distances[63]) && (distances[31] < distances[64]) && (distances[31] < distances[65]) && (distances[31] < distances[66]) && (distances[31] < distances[67]) && (distances[31] < distances[68]) && (distances[31] < distances[69]) && (distances[31] < distances[70]) && (distances[31] < distances[71]) && (distances[31] < distances[72]) && (distances[31] < distances[73]) && (distances[31] < distances[74]) && (distances[31] < distances[75]) && (distances[31] < distances[76]) && (distances[31] < distances[77]) && (distances[31] < distances[78]) && (distances[31] < distances[79]) && (distances[31] < distances[80]) && (distances[31] < distances[81]) && (distances[31] < distances[82]) && (distances[31] < distances[83]) && (distances[31] < distances[84]) && (distances[31] < distances[85]) && (distances[31] < distances[86]) && (distances[31] < distances[87]) && (distances[31] < distances[88]) && (distances[31] < distances[89])) begin
        dout <= 31;
      end else if((distances[32] < distances[33]) && (distances[32] < distances[34]) && (distances[32] < distances[35]) && (distances[32] < distances[36]) && (distances[32] < distances[37]) && (distances[32] < distances[38]) && (distances[32] < distances[39]) && (distances[32] < distances[40]) && (distances[32] < distances[41]) && (distances[32] < distances[42]) && (distances[32] < distances[43]) && (distances[32] < distances[44]) && (distances[32] < distances[45]) && (distances[32] < distances[46]) && (distances[32] < distances[47]) && (distances[32] < distances[48]) && (distances[32] < distances[49]) && (distances[32] < distances[50]) && (distances[32] < distances[51]) && (distances[32] < distances[52]) && (distances[32] < distances[53]) && (distances[32] < distances[54]) && (distances[32] < distances[55]) && (distances[32] < distances[56]) && (distances[32] < distances[57]) && (distances[32] < distances[58]) && (distances[32] < distances[59]) && (distances[32] < distances[60]) && (distances[32] < distances[61]) && (distances[32] < distances[62]) && (distances[32] < distances[63]) && (distances[32] < distances[64]) && (distances[32] < distances[65]) && (distances[32] < distances[66]) && (distances[32] < distances[67]) && (distances[32] < distances[68]) && (distances[32] < distances[69]) && (distances[32] < distances[70]) && (distances[32] < distances[71]) && (distances[32] < distances[72]) && (distances[32] < distances[73]) && (distances[32] < distances[74]) && (distances[32] < distances[75]) && (distances[32] < distances[76]) && (distances[32] < distances[77]) && (distances[32] < distances[78]) && (distances[32] < distances[79]) && (distances[32] < distances[80]) && (distances[32] < distances[81]) && (distances[32] < distances[82]) && (distances[32] < distances[83]) && (distances[32] < distances[84]) && (distances[32] < distances[85]) && (distances[32] < distances[86]) && (distances[32] < distances[87]) && (distances[32] < distances[88]) && (distances[32] < distances[89])) begin
        dout <= 32;
      end else if((distances[33] < distances[34]) && (distances[33] < distances[35]) && (distances[33] < distances[36]) && (distances[33] < distances[37]) && (distances[33] < distances[38]) && (distances[33] < distances[39]) && (distances[33] < distances[40]) && (distances[33] < distances[41]) && (distances[33] < distances[42]) && (distances[33] < distances[43]) && (distances[33] < distances[44]) && (distances[33] < distances[45]) && (distances[33] < distances[46]) && (distances[33] < distances[47]) && (distances[33] < distances[48]) && (distances[33] < distances[49]) && (distances[33] < distances[50]) && (distances[33] < distances[51]) && (distances[33] < distances[52]) && (distances[33] < distances[53]) && (distances[33] < distances[54]) && (distances[33] < distances[55]) && (distances[33] < distances[56]) && (distances[33] < distances[57]) && (distances[33] < distances[58]) && (distances[33] < distances[59]) && (distances[33] < distances[60]) && (distances[33] < distances[61]) && (distances[33] < distances[62]) && (distances[33] < distances[63]) && (distances[33] < distances[64]) && (distances[33] < distances[65]) && (distances[33] < distances[66]) && (distances[33] < distances[67]) && (distances[33] < distances[68]) && (distances[33] < distances[69]) && (distances[33] < distances[70]) && (distances[33] < distances[71]) && (distances[33] < distances[72]) && (distances[33] < distances[73]) && (distances[33] < distances[74]) && (distances[33] < distances[75]) && (distances[33] < distances[76]) && (distances[33] < distances[77]) && (distances[33] < distances[78]) && (distances[33] < distances[79]) && (distances[33] < distances[80]) && (distances[33] < distances[81]) && (distances[33] < distances[82]) && (distances[33] < distances[83]) && (distances[33] < distances[84]) && (distances[33] < distances[85]) && (distances[33] < distances[86]) && (distances[33] < distances[87]) && (distances[33] < distances[88]) && (distances[33] < distances[89])) begin
        dout <= 33;
      end else if((distances[34] < distances[35]) && (distances[34] < distances[36]) && (distances[34] < distances[37]) && (distances[34] < distances[38]) && (distances[34] < distances[39]) && (distances[34] < distances[40]) && (distances[34] < distances[41]) && (distances[34] < distances[42]) && (distances[34] < distances[43]) && (distances[34] < distances[44]) && (distances[34] < distances[45]) && (distances[34] < distances[46]) && (distances[34] < distances[47]) && (distances[34] < distances[48]) && (distances[34] < distances[49]) && (distances[34] < distances[50]) && (distances[34] < distances[51]) && (distances[34] < distances[52]) && (distances[34] < distances[53]) && (distances[34] < distances[54]) && (distances[34] < distances[55]) && (distances[34] < distances[56]) && (distances[34] < distances[57]) && (distances[34] < distances[58]) && (distances[34] < distances[59]) && (distances[34] < distances[60]) && (distances[34] < distances[61]) && (distances[34] < distances[62]) && (distances[34] < distances[63]) && (distances[34] < distances[64]) && (distances[34] < distances[65]) && (distances[34] < distances[66]) && (distances[34] < distances[67]) && (distances[34] < distances[68]) && (distances[34] < distances[69]) && (distances[34] < distances[70]) && (distances[34] < distances[71]) && (distances[34] < distances[72]) && (distances[34] < distances[73]) && (distances[34] < distances[74]) && (distances[34] < distances[75]) && (distances[34] < distances[76]) && (distances[34] < distances[77]) && (distances[34] < distances[78]) && (distances[34] < distances[79]) && (distances[34] < distances[80]) && (distances[34] < distances[81]) && (distances[34] < distances[82]) && (distances[34] < distances[83]) && (distances[34] < distances[84]) && (distances[34] < distances[85]) && (distances[34] < distances[86]) && (distances[34] < distances[87]) && (distances[34] < distances[88]) && (distances[34] < distances[89])) begin
        dout <= 34;
      end else if((distances[35] < distances[36]) && (distances[35] < distances[37]) && (distances[35] < distances[38]) && (distances[35] < distances[39]) && (distances[35] < distances[40]) && (distances[35] < distances[41]) && (distances[35] < distances[42]) && (distances[35] < distances[43]) && (distances[35] < distances[44]) && (distances[35] < distances[45]) && (distances[35] < distances[46]) && (distances[35] < distances[47]) && (distances[35] < distances[48]) && (distances[35] < distances[49]) && (distances[35] < distances[50]) && (distances[35] < distances[51]) && (distances[35] < distances[52]) && (distances[35] < distances[53]) && (distances[35] < distances[54]) && (distances[35] < distances[55]) && (distances[35] < distances[56]) && (distances[35] < distances[57]) && (distances[35] < distances[58]) && (distances[35] < distances[59]) && (distances[35] < distances[60]) && (distances[35] < distances[61]) && (distances[35] < distances[62]) && (distances[35] < distances[63]) && (distances[35] < distances[64]) && (distances[35] < distances[65]) && (distances[35] < distances[66]) && (distances[35] < distances[67]) && (distances[35] < distances[68]) && (distances[35] < distances[69]) && (distances[35] < distances[70]) && (distances[35] < distances[71]) && (distances[35] < distances[72]) && (distances[35] < distances[73]) && (distances[35] < distances[74]) && (distances[35] < distances[75]) && (distances[35] < distances[76]) && (distances[35] < distances[77]) && (distances[35] < distances[78]) && (distances[35] < distances[79]) && (distances[35] < distances[80]) && (distances[35] < distances[81]) && (distances[35] < distances[82]) && (distances[35] < distances[83]) && (distances[35] < distances[84]) && (distances[35] < distances[85]) && (distances[35] < distances[86]) && (distances[35] < distances[87]) && (distances[35] < distances[88]) && (distances[35] < distances[89])) begin
        dout <= 35;
      end else if((distances[36] < distances[37]) && (distances[36] < distances[38]) && (distances[36] < distances[39]) && (distances[36] < distances[40]) && (distances[36] < distances[41]) && (distances[36] < distances[42]) && (distances[36] < distances[43]) && (distances[36] < distances[44]) && (distances[36] < distances[45]) && (distances[36] < distances[46]) && (distances[36] < distances[47]) && (distances[36] < distances[48]) && (distances[36] < distances[49]) && (distances[36] < distances[50]) && (distances[36] < distances[51]) && (distances[36] < distances[52]) && (distances[36] < distances[53]) && (distances[36] < distances[54]) && (distances[36] < distances[55]) && (distances[36] < distances[56]) && (distances[36] < distances[57]) && (distances[36] < distances[58]) && (distances[36] < distances[59]) && (distances[36] < distances[60]) && (distances[36] < distances[61]) && (distances[36] < distances[62]) && (distances[36] < distances[63]) && (distances[36] < distances[64]) && (distances[36] < distances[65]) && (distances[36] < distances[66]) && (distances[36] < distances[67]) && (distances[36] < distances[68]) && (distances[36] < distances[69]) && (distances[36] < distances[70]) && (distances[36] < distances[71]) && (distances[36] < distances[72]) && (distances[36] < distances[73]) && (distances[36] < distances[74]) && (distances[36] < distances[75]) && (distances[36] < distances[76]) && (distances[36] < distances[77]) && (distances[36] < distances[78]) && (distances[36] < distances[79]) && (distances[36] < distances[80]) && (distances[36] < distances[81]) && (distances[36] < distances[82]) && (distances[36] < distances[83]) && (distances[36] < distances[84]) && (distances[36] < distances[85]) && (distances[36] < distances[86]) && (distances[36] < distances[87]) && (distances[36] < distances[88]) && (distances[36] < distances[89])) begin
        dout <= 36;
      end else if((distances[37] < distances[38]) && (distances[37] < distances[39]) && (distances[37] < distances[40]) && (distances[37] < distances[41]) && (distances[37] < distances[42]) && (distances[37] < distances[43]) && (distances[37] < distances[44]) && (distances[37] < distances[45]) && (distances[37] < distances[46]) && (distances[37] < distances[47]) && (distances[37] < distances[48]) && (distances[37] < distances[49]) && (distances[37] < distances[50]) && (distances[37] < distances[51]) && (distances[37] < distances[52]) && (distances[37] < distances[53]) && (distances[37] < distances[54]) && (distances[37] < distances[55]) && (distances[37] < distances[56]) && (distances[37] < distances[57]) && (distances[37] < distances[58]) && (distances[37] < distances[59]) && (distances[37] < distances[60]) && (distances[37] < distances[61]) && (distances[37] < distances[62]) && (distances[37] < distances[63]) && (distances[37] < distances[64]) && (distances[37] < distances[65]) && (distances[37] < distances[66]) && (distances[37] < distances[67]) && (distances[37] < distances[68]) && (distances[37] < distances[69]) && (distances[37] < distances[70]) && (distances[37] < distances[71]) && (distances[37] < distances[72]) && (distances[37] < distances[73]) && (distances[37] < distances[74]) && (distances[37] < distances[75]) && (distances[37] < distances[76]) && (distances[37] < distances[77]) && (distances[37] < distances[78]) && (distances[37] < distances[79]) && (distances[37] < distances[80]) && (distances[37] < distances[81]) && (distances[37] < distances[82]) && (distances[37] < distances[83]) && (distances[37] < distances[84]) && (distances[37] < distances[85]) && (distances[37] < distances[86]) && (distances[37] < distances[87]) && (distances[37] < distances[88]) && (distances[37] < distances[89])) begin
        dout <= 37;
      end else if((distances[38] < distances[39]) && (distances[38] < distances[40]) && (distances[38] < distances[41]) && (distances[38] < distances[42]) && (distances[38] < distances[43]) && (distances[38] < distances[44]) && (distances[38] < distances[45]) && (distances[38] < distances[46]) && (distances[38] < distances[47]) && (distances[38] < distances[48]) && (distances[38] < distances[49]) && (distances[38] < distances[50]) && (distances[38] < distances[51]) && (distances[38] < distances[52]) && (distances[38] < distances[53]) && (distances[38] < distances[54]) && (distances[38] < distances[55]) && (distances[38] < distances[56]) && (distances[38] < distances[57]) && (distances[38] < distances[58]) && (distances[38] < distances[59]) && (distances[38] < distances[60]) && (distances[38] < distances[61]) && (distances[38] < distances[62]) && (distances[38] < distances[63]) && (distances[38] < distances[64]) && (distances[38] < distances[65]) && (distances[38] < distances[66]) && (distances[38] < distances[67]) && (distances[38] < distances[68]) && (distances[38] < distances[69]) && (distances[38] < distances[70]) && (distances[38] < distances[71]) && (distances[38] < distances[72]) && (distances[38] < distances[73]) && (distances[38] < distances[74]) && (distances[38] < distances[75]) && (distances[38] < distances[76]) && (distances[38] < distances[77]) && (distances[38] < distances[78]) && (distances[38] < distances[79]) && (distances[38] < distances[80]) && (distances[38] < distances[81]) && (distances[38] < distances[82]) && (distances[38] < distances[83]) && (distances[38] < distances[84]) && (distances[38] < distances[85]) && (distances[38] < distances[86]) && (distances[38] < distances[87]) && (distances[38] < distances[88]) && (distances[38] < distances[89])) begin
        dout <= 38;
      end else if((distances[39] < distances[40]) && (distances[39] < distances[41]) && (distances[39] < distances[42]) && (distances[39] < distances[43]) && (distances[39] < distances[44]) && (distances[39] < distances[45]) && (distances[39] < distances[46]) && (distances[39] < distances[47]) && (distances[39] < distances[48]) && (distances[39] < distances[49]) && (distances[39] < distances[50]) && (distances[39] < distances[51]) && (distances[39] < distances[52]) && (distances[39] < distances[53]) && (distances[39] < distances[54]) && (distances[39] < distances[55]) && (distances[39] < distances[56]) && (distances[39] < distances[57]) && (distances[39] < distances[58]) && (distances[39] < distances[59]) && (distances[39] < distances[60]) && (distances[39] < distances[61]) && (distances[39] < distances[62]) && (distances[39] < distances[63]) && (distances[39] < distances[64]) && (distances[39] < distances[65]) && (distances[39] < distances[66]) && (distances[39] < distances[67]) && (distances[39] < distances[68]) && (distances[39] < distances[69]) && (distances[39] < distances[70]) && (distances[39] < distances[71]) && (distances[39] < distances[72]) && (distances[39] < distances[73]) && (distances[39] < distances[74]) && (distances[39] < distances[75]) && (distances[39] < distances[76]) && (distances[39] < distances[77]) && (distances[39] < distances[78]) && (distances[39] < distances[79]) && (distances[39] < distances[80]) && (distances[39] < distances[81]) && (distances[39] < distances[82]) && (distances[39] < distances[83]) && (distances[39] < distances[84]) && (distances[39] < distances[85]) && (distances[39] < distances[86]) && (distances[39] < distances[87]) && (distances[39] < distances[88]) && (distances[39] < distances[89])) begin
        dout <= 39;
      end else if((distances[40] < distances[41]) && (distances[40] < distances[42]) && (distances[40] < distances[43]) && (distances[40] < distances[44]) && (distances[40] < distances[45]) && (distances[40] < distances[46]) && (distances[40] < distances[47]) && (distances[40] < distances[48]) && (distances[40] < distances[49]) && (distances[40] < distances[50]) && (distances[40] < distances[51]) && (distances[40] < distances[52]) && (distances[40] < distances[53]) && (distances[40] < distances[54]) && (distances[40] < distances[55]) && (distances[40] < distances[56]) && (distances[40] < distances[57]) && (distances[40] < distances[58]) && (distances[40] < distances[59]) && (distances[40] < distances[60]) && (distances[40] < distances[61]) && (distances[40] < distances[62]) && (distances[40] < distances[63]) && (distances[40] < distances[64]) && (distances[40] < distances[65]) && (distances[40] < distances[66]) && (distances[40] < distances[67]) && (distances[40] < distances[68]) && (distances[40] < distances[69]) && (distances[40] < distances[70]) && (distances[40] < distances[71]) && (distances[40] < distances[72]) && (distances[40] < distances[73]) && (distances[40] < distances[74]) && (distances[40] < distances[75]) && (distances[40] < distances[76]) && (distances[40] < distances[77]) && (distances[40] < distances[78]) && (distances[40] < distances[79]) && (distances[40] < distances[80]) && (distances[40] < distances[81]) && (distances[40] < distances[82]) && (distances[40] < distances[83]) && (distances[40] < distances[84]) && (distances[40] < distances[85]) && (distances[40] < distances[86]) && (distances[40] < distances[87]) && (distances[40] < distances[88]) && (distances[40] < distances[89])) begin
        dout <= 40;
      end else if((distances[41] < distances[42]) && (distances[41] < distances[43]) && (distances[41] < distances[44]) && (distances[41] < distances[45]) && (distances[41] < distances[46]) && (distances[41] < distances[47]) && (distances[41] < distances[48]) && (distances[41] < distances[49]) && (distances[41] < distances[50]) && (distances[41] < distances[51]) && (distances[41] < distances[52]) && (distances[41] < distances[53]) && (distances[41] < distances[54]) && (distances[41] < distances[55]) && (distances[41] < distances[56]) && (distances[41] < distances[57]) && (distances[41] < distances[58]) && (distances[41] < distances[59]) && (distances[41] < distances[60]) && (distances[41] < distances[61]) && (distances[41] < distances[62]) && (distances[41] < distances[63]) && (distances[41] < distances[64]) && (distances[41] < distances[65]) && (distances[41] < distances[66]) && (distances[41] < distances[67]) && (distances[41] < distances[68]) && (distances[41] < distances[69]) && (distances[41] < distances[70]) && (distances[41] < distances[71]) && (distances[41] < distances[72]) && (distances[41] < distances[73]) && (distances[41] < distances[74]) && (distances[41] < distances[75]) && (distances[41] < distances[76]) && (distances[41] < distances[77]) && (distances[41] < distances[78]) && (distances[41] < distances[79]) && (distances[41] < distances[80]) && (distances[41] < distances[81]) && (distances[41] < distances[82]) && (distances[41] < distances[83]) && (distances[41] < distances[84]) && (distances[41] < distances[85]) && (distances[41] < distances[86]) && (distances[41] < distances[87]) && (distances[41] < distances[88]) && (distances[41] < distances[89])) begin
        dout <= 41;
      end else if((distances[42] < distances[43]) && (distances[42] < distances[44]) && (distances[42] < distances[45]) && (distances[42] < distances[46]) && (distances[42] < distances[47]) && (distances[42] < distances[48]) && (distances[42] < distances[49]) && (distances[42] < distances[50]) && (distances[42] < distances[51]) && (distances[42] < distances[52]) && (distances[42] < distances[53]) && (distances[42] < distances[54]) && (distances[42] < distances[55]) && (distances[42] < distances[56]) && (distances[42] < distances[57]) && (distances[42] < distances[58]) && (distances[42] < distances[59]) && (distances[42] < distances[60]) && (distances[42] < distances[61]) && (distances[42] < distances[62]) && (distances[42] < distances[63]) && (distances[42] < distances[64]) && (distances[42] < distances[65]) && (distances[42] < distances[66]) && (distances[42] < distances[67]) && (distances[42] < distances[68]) && (distances[42] < distances[69]) && (distances[42] < distances[70]) && (distances[42] < distances[71]) && (distances[42] < distances[72]) && (distances[42] < distances[73]) && (distances[42] < distances[74]) && (distances[42] < distances[75]) && (distances[42] < distances[76]) && (distances[42] < distances[77]) && (distances[42] < distances[78]) && (distances[42] < distances[79]) && (distances[42] < distances[80]) && (distances[42] < distances[81]) && (distances[42] < distances[82]) && (distances[42] < distances[83]) && (distances[42] < distances[84]) && (distances[42] < distances[85]) && (distances[42] < distances[86]) && (distances[42] < distances[87]) && (distances[42] < distances[88]) && (distances[42] < distances[89])) begin
        dout <= 42;
      end else if((distances[43] < distances[44]) && (distances[43] < distances[45]) && (distances[43] < distances[46]) && (distances[43] < distances[47]) && (distances[43] < distances[48]) && (distances[43] < distances[49]) && (distances[43] < distances[50]) && (distances[43] < distances[51]) && (distances[43] < distances[52]) && (distances[43] < distances[53]) && (distances[43] < distances[54]) && (distances[43] < distances[55]) && (distances[43] < distances[56]) && (distances[43] < distances[57]) && (distances[43] < distances[58]) && (distances[43] < distances[59]) && (distances[43] < distances[60]) && (distances[43] < distances[61]) && (distances[43] < distances[62]) && (distances[43] < distances[63]) && (distances[43] < distances[64]) && (distances[43] < distances[65]) && (distances[43] < distances[66]) && (distances[43] < distances[67]) && (distances[43] < distances[68]) && (distances[43] < distances[69]) && (distances[43] < distances[70]) && (distances[43] < distances[71]) && (distances[43] < distances[72]) && (distances[43] < distances[73]) && (distances[43] < distances[74]) && (distances[43] < distances[75]) && (distances[43] < distances[76]) && (distances[43] < distances[77]) && (distances[43] < distances[78]) && (distances[43] < distances[79]) && (distances[43] < distances[80]) && (distances[43] < distances[81]) && (distances[43] < distances[82]) && (distances[43] < distances[83]) && (distances[43] < distances[84]) && (distances[43] < distances[85]) && (distances[43] < distances[86]) && (distances[43] < distances[87]) && (distances[43] < distances[88]) && (distances[43] < distances[89])) begin
        dout <= 43;
      end else if((distances[44] < distances[45]) && (distances[44] < distances[46]) && (distances[44] < distances[47]) && (distances[44] < distances[48]) && (distances[44] < distances[49]) && (distances[44] < distances[50]) && (distances[44] < distances[51]) && (distances[44] < distances[52]) && (distances[44] < distances[53]) && (distances[44] < distances[54]) && (distances[44] < distances[55]) && (distances[44] < distances[56]) && (distances[44] < distances[57]) && (distances[44] < distances[58]) && (distances[44] < distances[59]) && (distances[44] < distances[60]) && (distances[44] < distances[61]) && (distances[44] < distances[62]) && (distances[44] < distances[63]) && (distances[44] < distances[64]) && (distances[44] < distances[65]) && (distances[44] < distances[66]) && (distances[44] < distances[67]) && (distances[44] < distances[68]) && (distances[44] < distances[69]) && (distances[44] < distances[70]) && (distances[44] < distances[71]) && (distances[44] < distances[72]) && (distances[44] < distances[73]) && (distances[44] < distances[74]) && (distances[44] < distances[75]) && (distances[44] < distances[76]) && (distances[44] < distances[77]) && (distances[44] < distances[78]) && (distances[44] < distances[79]) && (distances[44] < distances[80]) && (distances[44] < distances[81]) && (distances[44] < distances[82]) && (distances[44] < distances[83]) && (distances[44] < distances[84]) && (distances[44] < distances[85]) && (distances[44] < distances[86]) && (distances[44] < distances[87]) && (distances[44] < distances[88]) && (distances[44] < distances[89])) begin
        dout <= 44;
      end else if((distances[45] < distances[46]) && (distances[45] < distances[47]) && (distances[45] < distances[48]) && (distances[45] < distances[49]) && (distances[45] < distances[50]) && (distances[45] < distances[51]) && (distances[45] < distances[52]) && (distances[45] < distances[53]) && (distances[45] < distances[54]) && (distances[45] < distances[55]) && (distances[45] < distances[56]) && (distances[45] < distances[57]) && (distances[45] < distances[58]) && (distances[45] < distances[59]) && (distances[45] < distances[60]) && (distances[45] < distances[61]) && (distances[45] < distances[62]) && (distances[45] < distances[63]) && (distances[45] < distances[64]) && (distances[45] < distances[65]) && (distances[45] < distances[66]) && (distances[45] < distances[67]) && (distances[45] < distances[68]) && (distances[45] < distances[69]) && (distances[45] < distances[70]) && (distances[45] < distances[71]) && (distances[45] < distances[72]) && (distances[45] < distances[73]) && (distances[45] < distances[74]) && (distances[45] < distances[75]) && (distances[45] < distances[76]) && (distances[45] < distances[77]) && (distances[45] < distances[78]) && (distances[45] < distances[79]) && (distances[45] < distances[80]) && (distances[45] < distances[81]) && (distances[45] < distances[82]) && (distances[45] < distances[83]) && (distances[45] < distances[84]) && (distances[45] < distances[85]) && (distances[45] < distances[86]) && (distances[45] < distances[87]) && (distances[45] < distances[88]) && (distances[45] < distances[89])) begin
        dout <= 45;
      end else if((distances[46] < distances[47]) && (distances[46] < distances[48]) && (distances[46] < distances[49]) && (distances[46] < distances[50]) && (distances[46] < distances[51]) && (distances[46] < distances[52]) && (distances[46] < distances[53]) && (distances[46] < distances[54]) && (distances[46] < distances[55]) && (distances[46] < distances[56]) && (distances[46] < distances[57]) && (distances[46] < distances[58]) && (distances[46] < distances[59]) && (distances[46] < distances[60]) && (distances[46] < distances[61]) && (distances[46] < distances[62]) && (distances[46] < distances[63]) && (distances[46] < distances[64]) && (distances[46] < distances[65]) && (distances[46] < distances[66]) && (distances[46] < distances[67]) && (distances[46] < distances[68]) && (distances[46] < distances[69]) && (distances[46] < distances[70]) && (distances[46] < distances[71]) && (distances[46] < distances[72]) && (distances[46] < distances[73]) && (distances[46] < distances[74]) && (distances[46] < distances[75]) && (distances[46] < distances[76]) && (distances[46] < distances[77]) && (distances[46] < distances[78]) && (distances[46] < distances[79]) && (distances[46] < distances[80]) && (distances[46] < distances[81]) && (distances[46] < distances[82]) && (distances[46] < distances[83]) && (distances[46] < distances[84]) && (distances[46] < distances[85]) && (distances[46] < distances[86]) && (distances[46] < distances[87]) && (distances[46] < distances[88]) && (distances[46] < distances[89])) begin
        dout <= 46;
      end else if((distances[47] < distances[48]) && (distances[47] < distances[49]) && (distances[47] < distances[50]) && (distances[47] < distances[51]) && (distances[47] < distances[52]) && (distances[47] < distances[53]) && (distances[47] < distances[54]) && (distances[47] < distances[55]) && (distances[47] < distances[56]) && (distances[47] < distances[57]) && (distances[47] < distances[58]) && (distances[47] < distances[59]) && (distances[47] < distances[60]) && (distances[47] < distances[61]) && (distances[47] < distances[62]) && (distances[47] < distances[63]) && (distances[47] < distances[64]) && (distances[47] < distances[65]) && (distances[47] < distances[66]) && (distances[47] < distances[67]) && (distances[47] < distances[68]) && (distances[47] < distances[69]) && (distances[47] < distances[70]) && (distances[47] < distances[71]) && (distances[47] < distances[72]) && (distances[47] < distances[73]) && (distances[47] < distances[74]) && (distances[47] < distances[75]) && (distances[47] < distances[76]) && (distances[47] < distances[77]) && (distances[47] < distances[78]) && (distances[47] < distances[79]) && (distances[47] < distances[80]) && (distances[47] < distances[81]) && (distances[47] < distances[82]) && (distances[47] < distances[83]) && (distances[47] < distances[84]) && (distances[47] < distances[85]) && (distances[47] < distances[86]) && (distances[47] < distances[87]) && (distances[47] < distances[88]) && (distances[47] < distances[89])) begin
        dout <= 47;
      end else if((distances[48] < distances[49]) && (distances[48] < distances[50]) && (distances[48] < distances[51]) && (distances[48] < distances[52]) && (distances[48] < distances[53]) && (distances[48] < distances[54]) && (distances[48] < distances[55]) && (distances[48] < distances[56]) && (distances[48] < distances[57]) && (distances[48] < distances[58]) && (distances[48] < distances[59]) && (distances[48] < distances[60]) && (distances[48] < distances[61]) && (distances[48] < distances[62]) && (distances[48] < distances[63]) && (distances[48] < distances[64]) && (distances[48] < distances[65]) && (distances[48] < distances[66]) && (distances[48] < distances[67]) && (distances[48] < distances[68]) && (distances[48] < distances[69]) && (distances[48] < distances[70]) && (distances[48] < distances[71]) && (distances[48] < distances[72]) && (distances[48] < distances[73]) && (distances[48] < distances[74]) && (distances[48] < distances[75]) && (distances[48] < distances[76]) && (distances[48] < distances[77]) && (distances[48] < distances[78]) && (distances[48] < distances[79]) && (distances[48] < distances[80]) && (distances[48] < distances[81]) && (distances[48] < distances[82]) && (distances[48] < distances[83]) && (distances[48] < distances[84]) && (distances[48] < distances[85]) && (distances[48] < distances[86]) && (distances[48] < distances[87]) && (distances[48] < distances[88]) && (distances[48] < distances[89])) begin
        dout <= 48;
      end else if((distances[49] < distances[50]) && (distances[49] < distances[51]) && (distances[49] < distances[52]) && (distances[49] < distances[53]) && (distances[49] < distances[54]) && (distances[49] < distances[55]) && (distances[49] < distances[56]) && (distances[49] < distances[57]) && (distances[49] < distances[58]) && (distances[49] < distances[59]) && (distances[49] < distances[60]) && (distances[49] < distances[61]) && (distances[49] < distances[62]) && (distances[49] < distances[63]) && (distances[49] < distances[64]) && (distances[49] < distances[65]) && (distances[49] < distances[66]) && (distances[49] < distances[67]) && (distances[49] < distances[68]) && (distances[49] < distances[69]) && (distances[49] < distances[70]) && (distances[49] < distances[71]) && (distances[49] < distances[72]) && (distances[49] < distances[73]) && (distances[49] < distances[74]) && (distances[49] < distances[75]) && (distances[49] < distances[76]) && (distances[49] < distances[77]) && (distances[49] < distances[78]) && (distances[49] < distances[79]) && (distances[49] < distances[80]) && (distances[49] < distances[81]) && (distances[49] < distances[82]) && (distances[49] < distances[83]) && (distances[49] < distances[84]) && (distances[49] < distances[85]) && (distances[49] < distances[86]) && (distances[49] < distances[87]) && (distances[49] < distances[88]) && (distances[49] < distances[89])) begin
        dout <= 49;
      end else if((distances[50] < distances[51]) && (distances[50] < distances[52]) && (distances[50] < distances[53]) && (distances[50] < distances[54]) && (distances[50] < distances[55]) && (distances[50] < distances[56]) && (distances[50] < distances[57]) && (distances[50] < distances[58]) && (distances[50] < distances[59]) && (distances[50] < distances[60]) && (distances[50] < distances[61]) && (distances[50] < distances[62]) && (distances[50] < distances[63]) && (distances[50] < distances[64]) && (distances[50] < distances[65]) && (distances[50] < distances[66]) && (distances[50] < distances[67]) && (distances[50] < distances[68]) && (distances[50] < distances[69]) && (distances[50] < distances[70]) && (distances[50] < distances[71]) && (distances[50] < distances[72]) && (distances[50] < distances[73]) && (distances[50] < distances[74]) && (distances[50] < distances[75]) && (distances[50] < distances[76]) && (distances[50] < distances[77]) && (distances[50] < distances[78]) && (distances[50] < distances[79]) && (distances[50] < distances[80]) && (distances[50] < distances[81]) && (distances[50] < distances[82]) && (distances[50] < distances[83]) && (distances[50] < distances[84]) && (distances[50] < distances[85]) && (distances[50] < distances[86]) && (distances[50] < distances[87]) && (distances[50] < distances[88]) && (distances[50] < distances[89])) begin
        dout <= 50;
      end else if((distances[51] < distances[52]) && (distances[51] < distances[53]) && (distances[51] < distances[54]) && (distances[51] < distances[55]) && (distances[51] < distances[56]) && (distances[51] < distances[57]) && (distances[51] < distances[58]) && (distances[51] < distances[59]) && (distances[51] < distances[60]) && (distances[51] < distances[61]) && (distances[51] < distances[62]) && (distances[51] < distances[63]) && (distances[51] < distances[64]) && (distances[51] < distances[65]) && (distances[51] < distances[66]) && (distances[51] < distances[67]) && (distances[51] < distances[68]) && (distances[51] < distances[69]) && (distances[51] < distances[70]) && (distances[51] < distances[71]) && (distances[51] < distances[72]) && (distances[51] < distances[73]) && (distances[51] < distances[74]) && (distances[51] < distances[75]) && (distances[51] < distances[76]) && (distances[51] < distances[77]) && (distances[51] < distances[78]) && (distances[51] < distances[79]) && (distances[51] < distances[80]) && (distances[51] < distances[81]) && (distances[51] < distances[82]) && (distances[51] < distances[83]) && (distances[51] < distances[84]) && (distances[51] < distances[85]) && (distances[51] < distances[86]) && (distances[51] < distances[87]) && (distances[51] < distances[88]) && (distances[51] < distances[89])) begin
        dout <= 51;
      end else if((distances[52] < distances[53]) && (distances[52] < distances[54]) && (distances[52] < distances[55]) && (distances[52] < distances[56]) && (distances[52] < distances[57]) && (distances[52] < distances[58]) && (distances[52] < distances[59]) && (distances[52] < distances[60]) && (distances[52] < distances[61]) && (distances[52] < distances[62]) && (distances[52] < distances[63]) && (distances[52] < distances[64]) && (distances[52] < distances[65]) && (distances[52] < distances[66]) && (distances[52] < distances[67]) && (distances[52] < distances[68]) && (distances[52] < distances[69]) && (distances[52] < distances[70]) && (distances[52] < distances[71]) && (distances[52] < distances[72]) && (distances[52] < distances[73]) && (distances[52] < distances[74]) && (distances[52] < distances[75]) && (distances[52] < distances[76]) && (distances[52] < distances[77]) && (distances[52] < distances[78]) && (distances[52] < distances[79]) && (distances[52] < distances[80]) && (distances[52] < distances[81]) && (distances[52] < distances[82]) && (distances[52] < distances[83]) && (distances[52] < distances[84]) && (distances[52] < distances[85]) && (distances[52] < distances[86]) && (distances[52] < distances[87]) && (distances[52] < distances[88]) && (distances[52] < distances[89])) begin
        dout <= 52;
      end else if((distances[53] < distances[54]) && (distances[53] < distances[55]) && (distances[53] < distances[56]) && (distances[53] < distances[57]) && (distances[53] < distances[58]) && (distances[53] < distances[59]) && (distances[53] < distances[60]) && (distances[53] < distances[61]) && (distances[53] < distances[62]) && (distances[53] < distances[63]) && (distances[53] < distances[64]) && (distances[53] < distances[65]) && (distances[53] < distances[66]) && (distances[53] < distances[67]) && (distances[53] < distances[68]) && (distances[53] < distances[69]) && (distances[53] < distances[70]) && (distances[53] < distances[71]) && (distances[53] < distances[72]) && (distances[53] < distances[73]) && (distances[53] < distances[74]) && (distances[53] < distances[75]) && (distances[53] < distances[76]) && (distances[53] < distances[77]) && (distances[53] < distances[78]) && (distances[53] < distances[79]) && (distances[53] < distances[80]) && (distances[53] < distances[81]) && (distances[53] < distances[82]) && (distances[53] < distances[83]) && (distances[53] < distances[84]) && (distances[53] < distances[85]) && (distances[53] < distances[86]) && (distances[53] < distances[87]) && (distances[53] < distances[88]) && (distances[53] < distances[89])) begin
        dout <= 53;
      end else if((distances[54] < distances[55]) && (distances[54] < distances[56]) && (distances[54] < distances[57]) && (distances[54] < distances[58]) && (distances[54] < distances[59]) && (distances[54] < distances[60]) && (distances[54] < distances[61]) && (distances[54] < distances[62]) && (distances[54] < distances[63]) && (distances[54] < distances[64]) && (distances[54] < distances[65]) && (distances[54] < distances[66]) && (distances[54] < distances[67]) && (distances[54] < distances[68]) && (distances[54] < distances[69]) && (distances[54] < distances[70]) && (distances[54] < distances[71]) && (distances[54] < distances[72]) && (distances[54] < distances[73]) && (distances[54] < distances[74]) && (distances[54] < distances[75]) && (distances[54] < distances[76]) && (distances[54] < distances[77]) && (distances[54] < distances[78]) && (distances[54] < distances[79]) && (distances[54] < distances[80]) && (distances[54] < distances[81]) && (distances[54] < distances[82]) && (distances[54] < distances[83]) && (distances[54] < distances[84]) && (distances[54] < distances[85]) && (distances[54] < distances[86]) && (distances[54] < distances[87]) && (distances[54] < distances[88]) && (distances[54] < distances[89])) begin
        dout <= 54;
      end else if((distances[55] < distances[56]) && (distances[55] < distances[57]) && (distances[55] < distances[58]) && (distances[55] < distances[59]) && (distances[55] < distances[60]) && (distances[55] < distances[61]) && (distances[55] < distances[62]) && (distances[55] < distances[63]) && (distances[55] < distances[64]) && (distances[55] < distances[65]) && (distances[55] < distances[66]) && (distances[55] < distances[67]) && (distances[55] < distances[68]) && (distances[55] < distances[69]) && (distances[55] < distances[70]) && (distances[55] < distances[71]) && (distances[55] < distances[72]) && (distances[55] < distances[73]) && (distances[55] < distances[74]) && (distances[55] < distances[75]) && (distances[55] < distances[76]) && (distances[55] < distances[77]) && (distances[55] < distances[78]) && (distances[55] < distances[79]) && (distances[55] < distances[80]) && (distances[55] < distances[81]) && (distances[55] < distances[82]) && (distances[55] < distances[83]) && (distances[55] < distances[84]) && (distances[55] < distances[85]) && (distances[55] < distances[86]) && (distances[55] < distances[87]) && (distances[55] < distances[88]) && (distances[55] < distances[89])) begin
        dout <= 55;
      end else if((distances[56] < distances[57]) && (distances[56] < distances[58]) && (distances[56] < distances[59]) && (distances[56] < distances[60]) && (distances[56] < distances[61]) && (distances[56] < distances[62]) && (distances[56] < distances[63]) && (distances[56] < distances[64]) && (distances[56] < distances[65]) && (distances[56] < distances[66]) && (distances[56] < distances[67]) && (distances[56] < distances[68]) && (distances[56] < distances[69]) && (distances[56] < distances[70]) && (distances[56] < distances[71]) && (distances[56] < distances[72]) && (distances[56] < distances[73]) && (distances[56] < distances[74]) && (distances[56] < distances[75]) && (distances[56] < distances[76]) && (distances[56] < distances[77]) && (distances[56] < distances[78]) && (distances[56] < distances[79]) && (distances[56] < distances[80]) && (distances[56] < distances[81]) && (distances[56] < distances[82]) && (distances[56] < distances[83]) && (distances[56] < distances[84]) && (distances[56] < distances[85]) && (distances[56] < distances[86]) && (distances[56] < distances[87]) && (distances[56] < distances[88]) && (distances[56] < distances[89])) begin
        dout <= 56;
      end else if((distances[57] < distances[58]) && (distances[57] < distances[59]) && (distances[57] < distances[60]) && (distances[57] < distances[61]) && (distances[57] < distances[62]) && (distances[57] < distances[63]) && (distances[57] < distances[64]) && (distances[57] < distances[65]) && (distances[57] < distances[66]) && (distances[57] < distances[67]) && (distances[57] < distances[68]) && (distances[57] < distances[69]) && (distances[57] < distances[70]) && (distances[57] < distances[71]) && (distances[57] < distances[72]) && (distances[57] < distances[73]) && (distances[57] < distances[74]) && (distances[57] < distances[75]) && (distances[57] < distances[76]) && (distances[57] < distances[77]) && (distances[57] < distances[78]) && (distances[57] < distances[79]) && (distances[57] < distances[80]) && (distances[57] < distances[81]) && (distances[57] < distances[82]) && (distances[57] < distances[83]) && (distances[57] < distances[84]) && (distances[57] < distances[85]) && (distances[57] < distances[86]) && (distances[57] < distances[87]) && (distances[57] < distances[88]) && (distances[57] < distances[89])) begin
        dout <= 57;
      end else if((distances[58] < distances[59]) && (distances[58] < distances[60]) && (distances[58] < distances[61]) && (distances[58] < distances[62]) && (distances[58] < distances[63]) && (distances[58] < distances[64]) && (distances[58] < distances[65]) && (distances[58] < distances[66]) && (distances[58] < distances[67]) && (distances[58] < distances[68]) && (distances[58] < distances[69]) && (distances[58] < distances[70]) && (distances[58] < distances[71]) && (distances[58] < distances[72]) && (distances[58] < distances[73]) && (distances[58] < distances[74]) && (distances[58] < distances[75]) && (distances[58] < distances[76]) && (distances[58] < distances[77]) && (distances[58] < distances[78]) && (distances[58] < distances[79]) && (distances[58] < distances[80]) && (distances[58] < distances[81]) && (distances[58] < distances[82]) && (distances[58] < distances[83]) && (distances[58] < distances[84]) && (distances[58] < distances[85]) && (distances[58] < distances[86]) && (distances[58] < distances[87]) && (distances[58] < distances[88]) && (distances[58] < distances[89])) begin
        dout <= 58;
      end else if((distances[59] < distances[60]) && (distances[59] < distances[61]) && (distances[59] < distances[62]) && (distances[59] < distances[63]) && (distances[59] < distances[64]) && (distances[59] < distances[65]) && (distances[59] < distances[66]) && (distances[59] < distances[67]) && (distances[59] < distances[68]) && (distances[59] < distances[69]) && (distances[59] < distances[70]) && (distances[59] < distances[71]) && (distances[59] < distances[72]) && (distances[59] < distances[73]) && (distances[59] < distances[74]) && (distances[59] < distances[75]) && (distances[59] < distances[76]) && (distances[59] < distances[77]) && (distances[59] < distances[78]) && (distances[59] < distances[79]) && (distances[59] < distances[80]) && (distances[59] < distances[81]) && (distances[59] < distances[82]) && (distances[59] < distances[83]) && (distances[59] < distances[84]) && (distances[59] < distances[85]) && (distances[59] < distances[86]) && (distances[59] < distances[87]) && (distances[59] < distances[88]) && (distances[59] < distances[89])) begin
        dout <= 59;
      end else if((distances[60] < distances[61]) && (distances[60] < distances[62]) && (distances[60] < distances[63]) && (distances[60] < distances[64]) && (distances[60] < distances[65]) && (distances[60] < distances[66]) && (distances[60] < distances[67]) && (distances[60] < distances[68]) && (distances[60] < distances[69]) && (distances[60] < distances[70]) && (distances[60] < distances[71]) && (distances[60] < distances[72]) && (distances[60] < distances[73]) && (distances[60] < distances[74]) && (distances[60] < distances[75]) && (distances[60] < distances[76]) && (distances[60] < distances[77]) && (distances[60] < distances[78]) && (distances[60] < distances[79]) && (distances[60] < distances[80]) && (distances[60] < distances[81]) && (distances[60] < distances[82]) && (distances[60] < distances[83]) && (distances[60] < distances[84]) && (distances[60] < distances[85]) && (distances[60] < distances[86]) && (distances[60] < distances[87]) && (distances[60] < distances[88]) && (distances[60] < distances[89])) begin
        dout <= 60;
      end else if((distances[61] < distances[62]) && (distances[61] < distances[63]) && (distances[61] < distances[64]) && (distances[61] < distances[65]) && (distances[61] < distances[66]) && (distances[61] < distances[67]) && (distances[61] < distances[68]) && (distances[61] < distances[69]) && (distances[61] < distances[70]) && (distances[61] < distances[71]) && (distances[61] < distances[72]) && (distances[61] < distances[73]) && (distances[61] < distances[74]) && (distances[61] < distances[75]) && (distances[61] < distances[76]) && (distances[61] < distances[77]) && (distances[61] < distances[78]) && (distances[61] < distances[79]) && (distances[61] < distances[80]) && (distances[61] < distances[81]) && (distances[61] < distances[82]) && (distances[61] < distances[83]) && (distances[61] < distances[84]) && (distances[61] < distances[85]) && (distances[61] < distances[86]) && (distances[61] < distances[87]) && (distances[61] < distances[88]) && (distances[61] < distances[89])) begin
        dout <= 61;
      end else if((distances[62] < distances[63]) && (distances[62] < distances[64]) && (distances[62] < distances[65]) && (distances[62] < distances[66]) && (distances[62] < distances[67]) && (distances[62] < distances[68]) && (distances[62] < distances[69]) && (distances[62] < distances[70]) && (distances[62] < distances[71]) && (distances[62] < distances[72]) && (distances[62] < distances[73]) && (distances[62] < distances[74]) && (distances[62] < distances[75]) && (distances[62] < distances[76]) && (distances[62] < distances[77]) && (distances[62] < distances[78]) && (distances[62] < distances[79]) && (distances[62] < distances[80]) && (distances[62] < distances[81]) && (distances[62] < distances[82]) && (distances[62] < distances[83]) && (distances[62] < distances[84]) && (distances[62] < distances[85]) && (distances[62] < distances[86]) && (distances[62] < distances[87]) && (distances[62] < distances[88]) && (distances[62] < distances[89])) begin
        dout <= 62;
      end else if((distances[63] < distances[64]) && (distances[63] < distances[65]) && (distances[63] < distances[66]) && (distances[63] < distances[67]) && (distances[63] < distances[68]) && (distances[63] < distances[69]) && (distances[63] < distances[70]) && (distances[63] < distances[71]) && (distances[63] < distances[72]) && (distances[63] < distances[73]) && (distances[63] < distances[74]) && (distances[63] < distances[75]) && (distances[63] < distances[76]) && (distances[63] < distances[77]) && (distances[63] < distances[78]) && (distances[63] < distances[79]) && (distances[63] < distances[80]) && (distances[63] < distances[81]) && (distances[63] < distances[82]) && (distances[63] < distances[83]) && (distances[63] < distances[84]) && (distances[63] < distances[85]) && (distances[63] < distances[86]) && (distances[63] < distances[87]) && (distances[63] < distances[88]) && (distances[63] < distances[89])) begin
        dout <= 63;
      end else if((distances[64] < distances[65]) && (distances[64] < distances[66]) && (distances[64] < distances[67]) && (distances[64] < distances[68]) && (distances[64] < distances[69]) && (distances[64] < distances[70]) && (distances[64] < distances[71]) && (distances[64] < distances[72]) && (distances[64] < distances[73]) && (distances[64] < distances[74]) && (distances[64] < distances[75]) && (distances[64] < distances[76]) && (distances[64] < distances[77]) && (distances[64] < distances[78]) && (distances[64] < distances[79]) && (distances[64] < distances[80]) && (distances[64] < distances[81]) && (distances[64] < distances[82]) && (distances[64] < distances[83]) && (distances[64] < distances[84]) && (distances[64] < distances[85]) && (distances[64] < distances[86]) && (distances[64] < distances[87]) && (distances[64] < distances[88]) && (distances[64] < distances[89])) begin
        dout <= 64;
      end else if((distances[65] < distances[66]) && (distances[65] < distances[67]) && (distances[65] < distances[68]) && (distances[65] < distances[69]) && (distances[65] < distances[70]) && (distances[65] < distances[71]) && (distances[65] < distances[72]) && (distances[65] < distances[73]) && (distances[65] < distances[74]) && (distances[65] < distances[75]) && (distances[65] < distances[76]) && (distances[65] < distances[77]) && (distances[65] < distances[78]) && (distances[65] < distances[79]) && (distances[65] < distances[80]) && (distances[65] < distances[81]) && (distances[65] < distances[82]) && (distances[65] < distances[83]) && (distances[65] < distances[84]) && (distances[65] < distances[85]) && (distances[65] < distances[86]) && (distances[65] < distances[87]) && (distances[65] < distances[88]) && (distances[65] < distances[89])) begin
        dout <= 65;
      end else if((distances[66] < distances[67]) && (distances[66] < distances[68]) && (distances[66] < distances[69]) && (distances[66] < distances[70]) && (distances[66] < distances[71]) && (distances[66] < distances[72]) && (distances[66] < distances[73]) && (distances[66] < distances[74]) && (distances[66] < distances[75]) && (distances[66] < distances[76]) && (distances[66] < distances[77]) && (distances[66] < distances[78]) && (distances[66] < distances[79]) && (distances[66] < distances[80]) && (distances[66] < distances[81]) && (distances[66] < distances[82]) && (distances[66] < distances[83]) && (distances[66] < distances[84]) && (distances[66] < distances[85]) && (distances[66] < distances[86]) && (distances[66] < distances[87]) && (distances[66] < distances[88]) && (distances[66] < distances[89])) begin
        dout <= 66;
      end else if((distances[67] < distances[68]) && (distances[67] < distances[69]) && (distances[67] < distances[70]) && (distances[67] < distances[71]) && (distances[67] < distances[72]) && (distances[67] < distances[73]) && (distances[67] < distances[74]) && (distances[67] < distances[75]) && (distances[67] < distances[76]) && (distances[67] < distances[77]) && (distances[67] < distances[78]) && (distances[67] < distances[79]) && (distances[67] < distances[80]) && (distances[67] < distances[81]) && (distances[67] < distances[82]) && (distances[67] < distances[83]) && (distances[67] < distances[84]) && (distances[67] < distances[85]) && (distances[67] < distances[86]) && (distances[67] < distances[87]) && (distances[67] < distances[88]) && (distances[67] < distances[89])) begin
        dout <= 67;
      end else if((distances[68] < distances[69]) && (distances[68] < distances[70]) && (distances[68] < distances[71]) && (distances[68] < distances[72]) && (distances[68] < distances[73]) && (distances[68] < distances[74]) && (distances[68] < distances[75]) && (distances[68] < distances[76]) && (distances[68] < distances[77]) && (distances[68] < distances[78]) && (distances[68] < distances[79]) && (distances[68] < distances[80]) && (distances[68] < distances[81]) && (distances[68] < distances[82]) && (distances[68] < distances[83]) && (distances[68] < distances[84]) && (distances[68] < distances[85]) && (distances[68] < distances[86]) && (distances[68] < distances[87]) && (distances[68] < distances[88]) && (distances[68] < distances[89])) begin
        dout <= 68;
      end else if((distances[69] < distances[70]) && (distances[69] < distances[71]) && (distances[69] < distances[72]) && (distances[69] < distances[73]) && (distances[69] < distances[74]) && (distances[69] < distances[75]) && (distances[69] < distances[76]) && (distances[69] < distances[77]) && (distances[69] < distances[78]) && (distances[69] < distances[79]) && (distances[69] < distances[80]) && (distances[69] < distances[81]) && (distances[69] < distances[82]) && (distances[69] < distances[83]) && (distances[69] < distances[84]) && (distances[69] < distances[85]) && (distances[69] < distances[86]) && (distances[69] < distances[87]) && (distances[69] < distances[88]) && (distances[69] < distances[89])) begin
        dout <= 69;
      end else if((distances[70] < distances[71]) && (distances[70] < distances[72]) && (distances[70] < distances[73]) && (distances[70] < distances[74]) && (distances[70] < distances[75]) && (distances[70] < distances[76]) && (distances[70] < distances[77]) && (distances[70] < distances[78]) && (distances[70] < distances[79]) && (distances[70] < distances[80]) && (distances[70] < distances[81]) && (distances[70] < distances[82]) && (distances[70] < distances[83]) && (distances[70] < distances[84]) && (distances[70] < distances[85]) && (distances[70] < distances[86]) && (distances[70] < distances[87]) && (distances[70] < distances[88]) && (distances[70] < distances[89])) begin
        dout <= 70;
      end else if((distances[71] < distances[72]) && (distances[71] < distances[73]) && (distances[71] < distances[74]) && (distances[71] < distances[75]) && (distances[71] < distances[76]) && (distances[71] < distances[77]) && (distances[71] < distances[78]) && (distances[71] < distances[79]) && (distances[71] < distances[80]) && (distances[71] < distances[81]) && (distances[71] < distances[82]) && (distances[71] < distances[83]) && (distances[71] < distances[84]) && (distances[71] < distances[85]) && (distances[71] < distances[86]) && (distances[71] < distances[87]) && (distances[71] < distances[88]) && (distances[71] < distances[89])) begin
        dout <= 71;
      end else if((distances[72] < distances[73]) && (distances[72] < distances[74]) && (distances[72] < distances[75]) && (distances[72] < distances[76]) && (distances[72] < distances[77]) && (distances[72] < distances[78]) && (distances[72] < distances[79]) && (distances[72] < distances[80]) && (distances[72] < distances[81]) && (distances[72] < distances[82]) && (distances[72] < distances[83]) && (distances[72] < distances[84]) && (distances[72] < distances[85]) && (distances[72] < distances[86]) && (distances[72] < distances[87]) && (distances[72] < distances[88]) && (distances[72] < distances[89])) begin
        dout <= 72;
      end else if((distances[73] < distances[74]) && (distances[73] < distances[75]) && (distances[73] < distances[76]) && (distances[73] < distances[77]) && (distances[73] < distances[78]) && (distances[73] < distances[79]) && (distances[73] < distances[80]) && (distances[73] < distances[81]) && (distances[73] < distances[82]) && (distances[73] < distances[83]) && (distances[73] < distances[84]) && (distances[73] < distances[85]) && (distances[73] < distances[86]) && (distances[73] < distances[87]) && (distances[73] < distances[88]) && (distances[73] < distances[89])) begin
        dout <= 73;
      end else if((distances[74] < distances[75]) && (distances[74] < distances[76]) && (distances[74] < distances[77]) && (distances[74] < distances[78]) && (distances[74] < distances[79]) && (distances[74] < distances[80]) && (distances[74] < distances[81]) && (distances[74] < distances[82]) && (distances[74] < distances[83]) && (distances[74] < distances[84]) && (distances[74] < distances[85]) && (distances[74] < distances[86]) && (distances[74] < distances[87]) && (distances[74] < distances[88]) && (distances[74] < distances[89])) begin
        dout <= 74;
      end else if((distances[75] < distances[76]) && (distances[75] < distances[77]) && (distances[75] < distances[78]) && (distances[75] < distances[79]) && (distances[75] < distances[80]) && (distances[75] < distances[81]) && (distances[75] < distances[82]) && (distances[75] < distances[83]) && (distances[75] < distances[84]) && (distances[75] < distances[85]) && (distances[75] < distances[86]) && (distances[75] < distances[87]) && (distances[75] < distances[88]) && (distances[75] < distances[89])) begin
        dout <= 75;
      end else if((distances[76] < distances[77]) && (distances[76] < distances[78]) && (distances[76] < distances[79]) && (distances[76] < distances[80]) && (distances[76] < distances[81]) && (distances[76] < distances[82]) && (distances[76] < distances[83]) && (distances[76] < distances[84]) && (distances[76] < distances[85]) && (distances[76] < distances[86]) && (distances[76] < distances[87]) && (distances[76] < distances[88]) && (distances[76] < distances[89])) begin
        dout <= 76;
      end else if((distances[77] < distances[78]) && (distances[77] < distances[79]) && (distances[77] < distances[80]) && (distances[77] < distances[81]) && (distances[77] < distances[82]) && (distances[77] < distances[83]) && (distances[77] < distances[84]) && (distances[77] < distances[85]) && (distances[77] < distances[86]) && (distances[77] < distances[87]) && (distances[77] < distances[88]) && (distances[77] < distances[89])) begin
        dout <= 77;
      end else if((distances[78] < distances[79]) && (distances[78] < distances[80]) && (distances[78] < distances[81]) && (distances[78] < distances[82]) && (distances[78] < distances[83]) && (distances[78] < distances[84]) && (distances[78] < distances[85]) && (distances[78] < distances[86]) && (distances[78] < distances[87]) && (distances[78] < distances[88]) && (distances[78] < distances[89])) begin
        dout <= 78;
      end else if((distances[79] < distances[80]) && (distances[79] < distances[81]) && (distances[79] < distances[82]) && (distances[79] < distances[83]) && (distances[79] < distances[84]) && (distances[79] < distances[85]) && (distances[79] < distances[86]) && (distances[79] < distances[87]) && (distances[79] < distances[88]) && (distances[79] < distances[89])) begin
        dout <= 79;
      end else if((distances[80] < distances[81]) && (distances[80] < distances[82]) && (distances[80] < distances[83]) && (distances[80] < distances[84]) && (distances[80] < distances[85]) && (distances[80] < distances[86]) && (distances[80] < distances[87]) && (distances[80] < distances[88]) && (distances[80] < distances[89])) begin
        dout <= 80;
      end else if((distances[81] < distances[82]) && (distances[81] < distances[83]) && (distances[81] < distances[84]) && (distances[81] < distances[85]) && (distances[81] < distances[86]) && (distances[81] < distances[87]) && (distances[81] < distances[88]) && (distances[81] < distances[89])) begin
        dout <= 81;
      end else if((distances[82] < distances[83]) && (distances[82] < distances[84]) && (distances[82] < distances[85]) && (distances[82] < distances[86]) && (distances[82] < distances[87]) && (distances[82] < distances[88]) && (distances[82] < distances[89])) begin
        dout <= 82;
      end else if((distances[83] < distances[84]) && (distances[83] < distances[85]) && (distances[83] < distances[86]) && (distances[83] < distances[87]) && (distances[83] < distances[88]) && (distances[83] < distances[89])) begin
        dout <= 83;
      end else if((distances[84] < distances[85]) && (distances[84] < distances[86]) && (distances[84] < distances[87]) && (distances[84] < distances[88]) && (distances[84] < distances[89])) begin
        dout <= 84;
      end else if((distances[85] < distances[86]) && (distances[85] < distances[87]) && (distances[85] < distances[88]) && (distances[85] < distances[89])) begin
        dout <= 85;
      end else if((distances[86] < distances[87]) && (distances[86] < distances[88]) && (distances[86] < distances[89])) begin
        dout <= 86;
      end else if((distances[87] < distances[88]) && (distances[87] < distances[89])) begin
        dout <= 87;
      end else if((distances[88] < distances[89])) begin
        dout <= 88;
      end else if((distances[89] !=  distances[88])) begin
        dout <= 89;
      end else begin
        dout <= 90;
      end
    end
  end
endmodule