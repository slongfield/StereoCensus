/*  Basic population count for up to 128 bits. Could easily be extended to
 *  any power of two.
 * 
 *  Copyright (c) 2016, Stephen Longfield, stephenlongfield.com
 * 
 *  This program is free software: you can redistribute it and/or modify
 *  it under the terms of the GNU General Public License as published by
 *  the Free Software Foundation, either version 3 of the License, or
 *  (at your option) any later version.
 *
 *  This program is distributed in the hope that it will be useful,
 *  but WITHOUT ANY WARRANTY; without even the implied warranty of
 *  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *  GNU General Public License for more details.
 *
 *  You should have received a copy of the GNU General Public License
 *  along with this program.  If not, see <http://www.gnu.org/licenses/>.
 *
 */

`ifndef CENSUS_POP_COUNT_V_
`define CENSUS_POP_COUNT_V_

`timescale 1ns/1ps

`include "dff.v"

// pop_count computes the population count of the input.
module pop_count#(
  parameter WIDTH=1
  ) (
    input wire clk,
    input wire rst,

    input wire  [WIDTH-1:0] inp,
    output wire [WIDTH-1:0] outp
  );

  // Binary 010101010...
  localparam m1   = 128'h55555555555555555555555555555555;
  // Binary 0011001100...
  localparam m2   = 128'h33333333333333333333333333333333;
  // Binary 000011110000..
  localparam m4   = 128'h0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f;
  // Binary 0000000011111111...
  localparam m8   = 128'h00ff00ff00ff00ff00ff00ff00ff00ff;
  // And so on.
  localparam m16  = 128'h0000ffff0000ffff0000ffff0000ffff;
  localparam m32  = 128'h00000000ffffffff00000000ffffffff;
  localparam m64  = 128'h0000000000000000ffffffffffffffff;

  // Need to turn off of this lint check due to long-standing Veriloator bug#63.
  /* verilator lint_off UNOPTFLAT */
  wire [WIDTH-1:0] x[$clog2(WIDTH)];

  dff#(.WIDTH(WIDTH)) out_ff(clk, rst, x[$clog2(WIDTH)-1], outp);

  assign x[0] = (inp & m1[WIDTH-1:0]) + ((inp >> 1) & m1[WIDTH-1:0]);

  // This sequence of shifts and additions creates a simple unpipelined tree adder.
  // TODO(slongfield): Make this generated by a separate script.
  generate
  if ($clog2(WIDTH) >= 2) begin
    assign x[1] = (x[0] & m2[WIDTH-1:0]) + ((x[0] >> 2) & m2[WIDTH-1:0]);  
  end
  if ($clog2(WIDTH) >= 3) begin
    assign x[2] = (x[1] & m4[WIDTH-1:0]) + ((x[1] >> 4) & m4[WIDTH-1:0]);  
  end
  if ($clog2(WIDTH) >= 4) begin
    assign x[3] = (x[2] & m8[WIDTH-1:0]) + ((x[2] >> 8) & m8[WIDTH-1:0]);  
  end
  if ($clog2(WIDTH) >= 5) begin
    assign x[4] = (x[3] & m16[WIDTH-1:0]) + ((x[3] >> 16) & m16[WIDTH-1:0]);  
  end
  if ($clog2(WIDTH) >= 6) begin
    assign x[5] = (x[4] & m32[WIDTH-1:0]) + ((x[4] >> 32) & m32[WIDTH-1:0]);  
  end
  if ($clog2(WIDTH) >= 7) begin
    assign x[6] = (x[5] & m64[WIDTH-1:0]) + ((x[5] >> 64) & m64[WIDTH-1:0]);  
  end
  if ($clog2(WIDTH) > 7) begin
    initial begin
      assert(0); // Cannot handle widths larger than 128.
    end
  end
  endgenerate
  /* verilator lint_on UNOPTFLAT */
endmodule

`endif // CENSUS_POP_COUNT_V_
